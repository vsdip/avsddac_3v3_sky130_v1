* SPICE3 file created from 7bitdac_layout.ext - technology: sky130A

.option scale=10000u

X0 switch_layout_0/dd switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1 switch_layout_0/dd switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2 switch_layout_0/dinb d6 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X3 switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X4 x1_out_v switch_layout_0/dd out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X5 out_v switch_layout_0/dinb x1_out_v switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X6 x2_out_v switch_layout_0/dd out_v switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X7 out_v switch_layout_0/dinb x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X8 6bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X9 6bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X10 6bitdac_layout_0/switch_layout_0/dinb d5 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X11 6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X12 6bitdac_layout_0/x1_out_v 6bitdac_layout_0/switch_layout_0/dd x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X13 x1_out_v 6bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/x1_out_v 6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X14 6bitdac_layout_0/x2_out_v 6bitdac_layout_0/switch_layout_0/dd x1_out_v 6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X15 x1_out_v 6bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X16 6bitdac_layout_0/x1_vref5 6bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X17 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X18 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X19 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X20 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X21 6bitdac_layout_0/5bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X22 6bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X23 6bitdac_layout_0/5bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X24 6bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X25 6bitdac_layout_0/5bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X26 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X27 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X28 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X29 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X30 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X31 6bitdac_layout_0/5bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X32 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X33 6bitdac_layout_0/5bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X34 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X35 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X36 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X37 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X38 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X39 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X40 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X41 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X42 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X43 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X44 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X45 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X46 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X47 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X48 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X49 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X50 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X51 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X52 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X53 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X54 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X55 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X56 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X57 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X58 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X59 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X60 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X61 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X62 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X63 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X64 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X65 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X66 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X67 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X68 inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X69 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X70 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X71 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X72 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X73 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X74 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X75 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X76 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X77 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X78 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X79 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X80 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X81 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X82 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X83 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X84 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X85 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X86 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X87 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X88 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X89 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X90 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X91 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X92 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X93 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X94 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X95 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X96 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X97 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X98 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X99 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X100 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X101 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X102 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X103 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X104 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X105 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X106 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X107 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X108 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X109 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X110 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X111 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X112 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X113 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X114 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X115 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X116 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X117 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X118 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X119 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X120 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X121 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X122 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X123 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X124 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X125 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X126 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X127 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X128 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X129 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X130 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X131 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X132 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X133 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X134 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X135 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X136 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X137 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X138 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X139 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X140 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X141 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X142 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X143 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X144 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X145 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X146 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X147 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X148 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X149 6bitdac_layout_0/5bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X150 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X151 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X152 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X153 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X154 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X155 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X156 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X157 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X158 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X159 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X160 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X161 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X162 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X163 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X164 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X165 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X166 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X167 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X168 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X169 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X170 6bitdac_layout_0/5bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X171 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X172 6bitdac_layout_0/5bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X173 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X174 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X175 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X176 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X177 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X178 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X179 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X180 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X181 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X182 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X183 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X184 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X185 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X186 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X187 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X188 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X189 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X190 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X191 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X192 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X193 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X194 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X195 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X196 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X197 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X198 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X199 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X200 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X201 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X202 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X203 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X204 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X205 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X206 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X207 6bitdac_layout_0/5bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X208 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X209 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X210 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X211 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X212 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X213 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X214 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X215 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X216 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X217 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X218 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X219 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X220 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X221 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X222 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X223 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X224 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X225 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X226 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X227 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X228 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X229 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X230 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X231 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X232 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X233 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X234 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X235 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X236 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X237 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X238 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X239 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X240 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X241 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X242 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X243 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X244 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X245 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X246 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X247 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X248 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X249 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X250 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X251 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X252 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X253 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X254 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X255 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X256 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X257 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X258 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X259 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X260 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X261 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X262 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X263 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X264 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X265 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X266 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X267 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X268 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X269 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X270 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X271 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X272 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X273 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X274 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X275 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X276 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X277 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X278 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X279 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X280 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X281 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X282 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X283 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X284 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X285 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X286 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X287 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X288 6bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X289 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X290 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X291 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X292 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X293 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X294 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X295 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X296 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X297 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X298 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X299 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X300 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X301 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X302 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X303 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X304 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X305 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X306 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X307 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X308 6bitdac_layout_0/5bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X309 6bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X310 6bitdac_layout_0/5bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X311 6bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X312 6bitdac_layout_0/5bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X313 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X314 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X315 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X316 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X317 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X318 6bitdac_layout_0/5bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X319 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X320 6bitdac_layout_0/5bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X321 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X322 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X323 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X324 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X325 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X326 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X327 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X328 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X329 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X330 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X331 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X332 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X333 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X334 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X335 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X336 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X337 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X338 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X339 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X340 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X341 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X342 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X343 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X344 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X345 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X346 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X347 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X348 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X349 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X350 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X351 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X352 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X353 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X354 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X355 6bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X356 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X357 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X358 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X359 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X360 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X361 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X362 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X363 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X364 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X365 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X366 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X367 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X368 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X369 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X370 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X371 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X372 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X373 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X374 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X375 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X376 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X377 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X378 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X379 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X380 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X381 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X382 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X383 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X384 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X385 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X386 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X387 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X388 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X389 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X390 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X391 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X392 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X393 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X394 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X395 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X396 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X397 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X398 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X399 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X400 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X401 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X402 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X403 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X404 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X405 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X406 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X407 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X408 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X409 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X410 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X411 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X412 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X413 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X414 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X415 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X416 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X417 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X418 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X419 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X420 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X421 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X422 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X423 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X424 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X425 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X426 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X427 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X428 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X429 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X430 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X431 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X432 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X433 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X434 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X435 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X436 6bitdac_layout_0/5bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X437 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X438 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X439 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X440 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X441 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X442 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X443 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X444 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X445 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X446 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X447 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X448 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X449 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X450 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X451 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X452 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X453 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X454 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X455 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X456 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X457 6bitdac_layout_0/5bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X458 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X459 6bitdac_layout_0/5bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X460 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X461 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X462 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X463 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X464 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X465 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X466 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X467 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X468 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X469 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X470 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X471 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X472 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X473 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X474 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X475 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X476 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X477 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X478 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X479 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X480 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X481 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X482 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X483 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X484 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X485 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X486 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X487 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X488 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X489 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X490 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X491 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X492 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X493 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X494 6bitdac_layout_0/5bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X495 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X496 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X497 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X498 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X499 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X500 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X501 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X502 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X503 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X504 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X505 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X506 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X507 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X508 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X509 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X510 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X511 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X512 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X513 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X514 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X515 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X516 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X517 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X518 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X519 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X520 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X521 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X522 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X523 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X524 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X525 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X526 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X527 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X528 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X529 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X530 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X531 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X532 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X533 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X534 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X535 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X536 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X537 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X538 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X539 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X540 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X541 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X542 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X543 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X544 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X545 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X546 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X547 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X548 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X549 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X550 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X551 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X552 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X553 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X554 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X555 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X556 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X557 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X558 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X559 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X560 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X561 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X562 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X563 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X564 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X565 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X566 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X567 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X568 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X569 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X570 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X571 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X572 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X573 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X574 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X575 x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X576 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X577 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X578 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X579 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X580 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X581 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X582 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X583 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X584 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X585 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X586 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X587 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X588 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X589 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X590 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X591 6bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X592 6bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X593 6bitdac_layout_1/switch_layout_0/dinb d5 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X594 6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X595 6bitdac_layout_1/x1_out_v 6bitdac_layout_1/switch_layout_0/dd x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X596 x2_out_v 6bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/x1_out_v 6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X597 6bitdac_layout_1/x2_out_v 6bitdac_layout_1/switch_layout_0/dd x2_out_v 6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X598 x2_out_v 6bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X599 6bitdac_layout_1/x1_vref5 6bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X600 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X601 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X602 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X603 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X604 6bitdac_layout_1/5bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X605 6bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X606 6bitdac_layout_1/5bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X607 6bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X608 6bitdac_layout_1/5bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X609 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X610 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X611 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X612 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X613 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X614 6bitdac_layout_1/5bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X615 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X616 6bitdac_layout_1/5bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X617 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X618 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X619 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X620 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X621 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X622 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X623 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X624 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X625 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X626 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X627 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X628 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X629 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X630 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X631 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X632 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X633 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X634 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X635 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X636 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X637 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X638 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X639 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X640 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X641 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X642 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X643 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X644 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X645 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X646 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X647 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X648 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X649 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X650 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X651 x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X652 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X653 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X654 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X655 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X656 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X657 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X658 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X659 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X660 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X661 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X662 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X663 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X664 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X665 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X666 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X667 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X668 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X669 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X670 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X671 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X672 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X673 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X674 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X675 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X676 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X677 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X678 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X679 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X680 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X681 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X682 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X683 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X684 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X685 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X686 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X687 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X688 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X689 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X690 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X691 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X692 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X693 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X694 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X695 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X696 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X697 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X698 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X699 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X700 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X701 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X702 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X703 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X704 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X705 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X706 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X707 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X708 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X709 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X710 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X711 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X712 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X713 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X714 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X715 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X716 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X717 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X718 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X719 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X720 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X721 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X722 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X723 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X724 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X725 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X726 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X727 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X728 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X729 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X730 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X731 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X732 6bitdac_layout_1/5bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X733 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X734 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X735 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X736 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X737 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X738 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X739 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X740 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X741 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X742 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X743 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X744 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X745 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X746 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X747 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X748 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X749 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X750 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X751 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X752 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X753 6bitdac_layout_1/5bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X754 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X755 6bitdac_layout_1/5bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X756 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X757 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X758 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X759 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X760 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X761 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X762 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X763 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X764 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X765 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X766 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X767 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X768 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X769 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X770 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X771 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X772 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X773 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X774 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X775 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X776 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X777 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X778 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X779 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X780 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X781 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X782 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X783 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X784 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X785 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X786 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X787 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X788 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X789 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X790 6bitdac_layout_1/5bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X791 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X792 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X793 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X794 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X795 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X796 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X797 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X798 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X799 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X800 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X801 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X802 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X803 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X804 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X805 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X806 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X807 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X808 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X809 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X810 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X811 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X812 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X813 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X814 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X815 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X816 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X817 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X818 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X819 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X820 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X821 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X822 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X823 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X824 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X825 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X826 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X827 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X828 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X829 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X830 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X831 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X832 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X833 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X834 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X835 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X836 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X837 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X838 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X839 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X840 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X841 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X842 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X843 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X844 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X845 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X846 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X847 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X848 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X849 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X850 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X851 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X852 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X853 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X854 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X855 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X856 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X857 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X858 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X859 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X860 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X861 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X862 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X863 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X864 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X865 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X866 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X867 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X868 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X869 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X870 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X871 6bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X872 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X873 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X874 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X875 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X876 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X877 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X878 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X879 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X880 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X881 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X882 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X883 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X884 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X885 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X886 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X887 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X888 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X889 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X890 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X891 6bitdac_layout_1/5bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X892 6bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X893 6bitdac_layout_1/5bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X894 6bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X895 6bitdac_layout_1/5bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X896 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X897 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X898 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X899 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X900 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X901 6bitdac_layout_1/5bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X902 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X903 6bitdac_layout_1/5bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X904 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X905 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X906 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X907 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X908 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X909 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X910 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X911 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X912 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X913 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X914 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X915 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X916 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X917 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X918 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X919 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X920 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X921 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X922 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X923 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X924 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X925 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X926 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X927 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X928 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X929 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X930 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X931 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X932 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X933 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X934 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X935 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X936 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X937 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X938 6bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X939 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X940 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X941 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X942 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X943 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X944 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X945 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X946 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X947 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X948 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X949 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X950 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X951 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X952 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X953 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X954 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X955 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X956 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X957 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X958 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X959 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X960 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X961 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X962 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X963 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X964 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X965 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X966 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X967 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X968 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X969 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X970 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X971 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X972 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X973 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X974 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X975 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X976 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X977 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X978 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X979 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X980 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X981 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X982 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X983 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X984 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X985 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X986 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X987 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X988 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X989 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X990 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X991 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X992 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X993 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X994 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X995 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X996 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X997 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X998 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X999 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1000 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1001 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1002 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1003 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1004 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1005 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1006 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1007 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1008 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1009 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1010 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1011 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1012 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1013 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1014 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1015 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1016 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1017 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1018 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1019 6bitdac_layout_1/5bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1020 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1021 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1022 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1023 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1024 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1025 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1026 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1027 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1028 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1029 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1030 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1031 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1032 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1033 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1034 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1035 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1036 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1037 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1038 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1039 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1040 6bitdac_layout_1/5bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1041 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1042 6bitdac_layout_1/5bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1043 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1044 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1045 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1046 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1047 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1048 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1049 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1050 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1051 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1052 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1053 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1054 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1055 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1056 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1057 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1058 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1059 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1060 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1061 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1062 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1063 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1064 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1065 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1066 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1067 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1068 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1069 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1070 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1071 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1072 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1073 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1074 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1075 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1076 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1077 6bitdac_layout_1/5bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1078 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1079 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1080 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1081 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1082 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1083 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1084 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1085 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1086 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1087 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1088 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1089 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1090 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1091 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1092 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1093 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1094 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1095 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1096 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1097 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1098 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1099 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1100 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1101 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1102 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1103 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1104 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1105 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1106 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1107 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1108 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1109 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1110 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1111 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1112 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1113 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1114 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1115 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1116 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1117 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1118 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1119 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1120 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1121 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1122 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1123 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1124 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1125 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1126 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1127 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1128 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1129 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1130 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1131 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1132 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1133 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1134 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1135 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1136 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1137 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1138 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1139 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1140 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1141 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1142 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1143 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1144 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1145 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1146 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1147 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1148 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1149 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1150 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1151 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1152 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1153 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1154 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1155 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1156 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1157 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1158 inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1159 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1160 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1161 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1162 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1163 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1164 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1165 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1166 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1167 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1168 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1169 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1170 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1171 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 inp2 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1172 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1173 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1174 x1_vref5 x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
C0 d5 d4 2.45fF
C1 d1 d0 11.80fF
C2 d1 d2 4.05fF
C3 vdd d0 6.67fF
C4 d4 d3 4.45fF
C5 vdd d2 2.22fF
C6 d2 d3 5.82fF
C7 d1 vdd 5.33fF
C8 vdd gnd 245.37fF
C9 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C10 6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C11 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C12 6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C13 x1_vref5 gnd 2.08fF
C14 d0 gnd 105.21fF
C15 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C16 6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C17 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C18 6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C19 d5 gnd 48.76fF
