magic
tech sky130A
timestamp 1616619357
<< locali >>
rect 9958 24341 9981 24343
rect 9958 24340 9982 24341
rect 9958 24337 9983 24340
rect 9958 24318 9962 24337
rect 9979 24335 9983 24337
rect 21880 24335 22581 24339
rect 9979 24320 22581 24335
rect 9979 24318 21919 24320
rect 9958 24316 21919 24318
rect 9958 24315 13627 24316
rect 22558 24312 22581 24320
rect 5884 24048 10081 24050
rect -126 24025 10430 24048
rect -126 24023 5909 24025
rect -126 24020 1724 24023
rect -123 -82 -97 24020
rect 272 23923 301 24003
rect 9958 23992 9988 23995
rect 9958 23973 9965 23992
rect 9982 23973 9988 23992
rect 9958 23970 9988 23973
rect 9959 15390 9982 23970
rect 10405 23910 10429 24025
rect 22558 23070 22583 24312
rect 9959 15372 9985 15390
rect 9961 13692 9985 15372
rect 9958 13671 9985 13692
rect 9958 13348 9982 13671
rect 9958 13331 9983 13348
rect 9959 13002 9983 13331
rect 22558 13120 22585 23070
rect 22558 13102 22590 13120
rect 9959 12987 9985 13002
rect 9961 12293 9985 12987
rect 22560 12852 22590 13102
rect 22561 12675 22588 12852
rect 22658 12535 22781 12543
rect 22658 12513 22668 12535
rect 22689 12513 22781 12535
rect 22658 12509 22781 12513
rect 21442 12424 21484 12476
rect 20802 12305 21185 12307
rect 20089 12277 21186 12305
rect 20089 12275 20847 12277
rect 8630 6736 8690 12258
rect 8630 6699 8642 6736
rect 8675 6699 8690 6736
rect 8630 6690 8690 6699
rect 18798 6675 18819 12242
rect 21166 12081 21186 12277
rect 22588 12083 22608 12301
rect 21942 12081 22611 12083
rect 21166 12061 22611 12081
rect 21166 12060 22346 12061
rect 21166 12058 21962 12060
rect 18798 6652 18801 6675
rect 18818 6652 18819 6675
rect 18798 6647 18819 6652
rect 6968 6498 7022 6552
rect 8615 6517 8680 6523
rect 6973 4645 7017 6498
rect 8615 6480 8632 6517
rect 8665 6480 8680 6517
rect 8615 5851 8680 6480
rect 8615 5757 8684 5851
rect 6964 4065 7017 4645
rect 6964 3730 7008 4065
rect 6964 3410 7012 3730
rect 6964 3388 6979 3410
rect 6965 3383 6979 3388
rect 7000 3383 7012 3410
rect 6965 3370 7012 3383
rect 5417 3142 5559 3191
rect 5419 2725 5454 3142
rect 5415 2692 5454 2725
rect 6964 3113 7008 3139
rect 6964 3086 6974 3113
rect 6995 3086 7008 3113
rect 5415 2388 5452 2692
rect 5412 2237 5452 2388
rect 5412 1937 5449 2237
rect 6964 2062 7008 3086
rect 6965 2026 7006 2062
rect 6965 1959 7021 2026
rect 5412 1913 5421 1937
rect 5441 1913 5449 1937
rect 5412 1900 5449 1913
rect 3742 1734 3791 1776
rect 5406 1769 5443 1780
rect 5406 1745 5408 1769
rect 5428 1745 5443 1769
rect 3743 1456 3770 1734
rect 3741 1063 3771 1456
rect 5406 1437 5443 1745
rect 3741 1035 3746 1063
rect 3764 1035 3771 1063
rect 3741 1015 3771 1035
rect 3741 875 3771 880
rect 1991 853 2004 862
rect 1991 602 2020 853
rect 1991 583 1995 602
rect 2017 583 2020 602
rect 1991 577 2020 583
rect 3741 847 3746 875
rect 3764 847 3771 875
rect 3741 537 3771 847
rect 1985 507 2022 511
rect 471 477 515 490
rect 1985 488 1993 507
rect 2015 488 2022 507
rect 471 350 506 477
rect 1985 465 2022 488
rect 3734 500 3771 537
rect 1985 398 2020 465
rect 471 346 505 350
rect 472 317 505 346
rect 1983 345 2020 398
rect 472 302 504 317
rect 468 299 504 302
rect 1983 300 2010 345
rect 468 280 474 299
rect 496 280 504 299
rect 468 275 504 280
rect 472 206 506 209
rect 472 204 509 206
rect 472 185 479 204
rect 501 185 509 204
rect 472 182 509 185
rect 472 179 505 182
rect 474 145 505 179
rect 474 84 506 145
rect 21 -1 107 17
rect 21 -59 52 -1
rect 472 -14 506 84
rect 1969 38 2010 300
rect 3734 196 3769 500
rect 5405 197 5449 1437
rect 6967 569 7021 1959
rect 8624 695 8684 5757
rect 17122 3712 17144 6568
rect 18795 6468 18817 6481
rect 18795 6445 18798 6468
rect 18815 6445 18817 6468
rect 18795 6440 18817 6445
rect 17118 3655 17144 3712
rect 17118 3315 17143 3655
rect 17118 3295 17121 3315
rect 17138 3295 17143 3315
rect 17118 3289 17143 3295
rect 15504 3134 15693 3196
rect 15504 3080 15566 3134
rect 17121 3115 17143 3119
rect 17119 3114 17143 3115
rect 17119 3093 17121 3114
rect 17138 3093 17143 3114
rect 17119 3086 17143 3093
rect 15509 2013 15565 3080
rect 15501 1925 15572 2013
rect 15501 1892 15529 1925
rect 15552 1892 15572 1925
rect 15501 1867 15572 1892
rect 13888 1051 13927 1757
rect 13888 1016 13897 1051
rect 13923 1016 13927 1051
rect 13888 992 13927 1016
rect 15520 1709 15564 1724
rect 15520 1676 15532 1709
rect 15555 1676 15564 1709
rect 1969 19 2009 38
rect -123 -180 -96 -82
rect -123 -181 86 -180
rect 107 -181 154 -175
rect -123 -208 154 -181
rect -59 -209 154 -208
rect 107 -210 154 -209
rect 468 -784 506 -14
rect 468 -970 507 -784
rect 468 -1198 508 -970
rect 1965 -1012 2009 19
rect 3718 -975 3774 196
rect 5402 -894 5449 197
rect 6945 382 7021 569
rect 6945 -742 7006 382
rect 8614 -521 8704 695
rect 12125 626 12168 877
rect 12125 596 12138 626
rect 12161 596 12168 626
rect 12125 589 12168 596
rect 13883 815 13922 838
rect 13883 780 13888 815
rect 13914 780 13922 815
rect 12119 464 12162 492
rect 10599 288 10632 460
rect 10599 264 10603 288
rect 10621 264 10632 288
rect 12119 434 12132 464
rect 12155 434 12162 464
rect 10595 183 10628 187
rect 10595 158 10603 183
rect 10621 158 10628 183
rect 10595 34 10628 158
rect 10595 -9 10629 34
rect 10207 -64 10234 -14
rect 10606 -476 10629 -9
rect 12119 -30 12162 434
rect 13883 136 13922 780
rect 15520 766 15564 1676
rect 15516 483 15573 766
rect 15516 258 15588 483
rect 13856 73 13922 136
rect 12119 -456 12149 -30
rect 12118 -460 12149 -456
rect 10603 -483 10634 -476
rect 10603 -500 10608 -483
rect 10625 -500 10634 -483
rect 12118 -486 12124 -460
rect 12145 -486 12149 -460
rect 13856 -440 13905 73
rect 13856 -469 13862 -440
rect 13888 -469 13905 -440
rect 13856 -481 13905 -469
rect 15524 -415 15588 258
rect 17121 236 17143 3086
rect 18796 1056 18817 6440
rect 17101 209 17143 236
rect 17101 167 17148 209
rect 17105 -109 17148 167
rect 15524 -457 15540 -415
rect 15578 -457 15588 -415
rect 12118 -498 12149 -486
rect 15524 -489 15588 -457
rect 17101 -159 17148 -109
rect 17101 -449 17144 -159
rect 17101 -470 17107 -449
rect 17130 -470 17144 -449
rect 17101 -477 17144 -470
rect 10603 -503 10634 -500
rect 18766 -521 18826 1056
rect 8599 -600 18827 -521
rect 8599 -608 9549 -600
rect 13798 -611 18827 -600
rect 13798 -626 15973 -611
rect 16809 -735 17137 -726
rect 10208 -741 17137 -735
rect 10208 -742 17109 -741
rect 6945 -762 17109 -742
rect 17132 -762 17137 -741
rect 6945 -803 17137 -762
rect 6945 -810 10291 -803
rect 16809 -810 17137 -803
rect 14092 -870 15586 -863
rect 10622 -871 15586 -870
rect 10622 -878 15530 -871
rect 7185 -894 15530 -878
rect 5402 -913 15530 -894
rect 15568 -913 15586 -871
rect 5402 -927 15586 -913
rect 5402 -934 14204 -927
rect 5402 -942 10703 -934
rect 5402 -954 7209 -942
rect 5446 -958 7209 -954
rect 3706 -993 3776 -975
rect 5678 -992 5849 -988
rect 5678 -993 12289 -992
rect 3706 -1010 12289 -993
rect 1965 -1136 2005 -1012
rect 3706 -1020 13909 -1010
rect 3706 -1049 13870 -1020
rect 13896 -1049 13909 -1020
rect 3706 -1060 13909 -1049
rect 3706 -1062 12289 -1060
rect 3706 -1065 5750 -1062
rect 3706 -1074 3776 -1065
rect 1964 -1138 2024 -1136
rect 6133 -1138 10382 -1130
rect 1964 -1164 12125 -1138
rect 12146 -1164 12150 -1138
rect 1964 -1171 12150 -1164
rect 1964 -1179 6199 -1171
rect 471 -1199 508 -1198
rect 10600 -1199 10630 -1195
rect 471 -1200 2043 -1199
rect 9802 -1200 10630 -1199
rect 471 -1202 10630 -1200
rect 471 -1220 10605 -1202
rect 10623 -1220 10630 -1202
rect 471 -1224 10630 -1220
rect 471 -1227 9871 -1224
rect 10600 -1226 10630 -1224
rect 471 -1228 508 -1227
rect 2030 -1228 9871 -1227
<< viali >>
rect 9962 24318 9979 24337
rect 9965 23973 9982 23992
rect 22668 12513 22689 12535
rect 8642 6699 8675 6736
rect 18801 6652 18818 6675
rect 8632 6480 8665 6517
rect 6979 3383 7000 3410
rect 6974 3086 6995 3113
rect 5421 1913 5441 1937
rect 5408 1745 5428 1769
rect 3746 1035 3764 1063
rect 1995 583 2017 602
rect 3746 847 3764 875
rect 1993 488 2015 507
rect 474 280 496 299
rect 479 185 501 204
rect 18798 6445 18815 6468
rect 17121 3295 17138 3315
rect 17121 3093 17138 3114
rect 15529 1892 15552 1925
rect 13897 1016 13923 1051
rect 15532 1676 15555 1709
rect 12138 596 12161 626
rect 13888 780 13914 815
rect 10603 263 10621 288
rect 12132 434 12155 464
rect 10603 158 10621 183
rect 10608 -500 10625 -483
rect 12124 -486 12145 -460
rect 13862 -469 13888 -440
rect 15540 -457 15578 -415
rect 17107 -470 17130 -449
rect 17109 -762 17132 -741
rect 15530 -913 15568 -871
rect 13870 -1049 13896 -1020
rect 12125 -1164 12146 -1138
rect 10605 -1220 10623 -1202
<< metal1 >>
rect 9958 24340 9981 24343
rect 9958 24337 9983 24340
rect 9958 24318 9962 24337
rect 9979 24318 9983 24337
rect 9958 24315 9983 24318
rect 9958 23995 9981 24315
rect 9958 23992 9988 23995
rect 9958 23973 9965 23992
rect 9982 23973 9988 23992
rect 9958 23970 9988 23973
rect 21887 12690 21941 12696
rect 21887 12662 21904 12690
rect 21933 12662 21941 12690
rect 21887 12658 21941 12662
rect 22658 12535 22696 12542
rect 22658 12513 22668 12535
rect 22689 12513 22696 12535
rect 22658 12509 22696 12513
rect 21525 12306 21567 12331
rect 21525 12276 21530 12306
rect 21559 12276 21567 12306
rect 21525 12259 21567 12276
rect 8615 6736 8689 6746
rect 8615 6699 8642 6736
rect 8675 6699 8689 6736
rect 8615 6517 8689 6699
rect 8615 6480 8632 6517
rect 8665 6480 8689 6517
rect 8615 6467 8689 6480
rect 18795 6675 18821 6682
rect 18795 6652 18801 6675
rect 18818 6652 18821 6675
rect 18795 6468 18821 6652
rect 18795 6445 18798 6468
rect 18815 6445 18821 6468
rect 18795 6439 18821 6445
rect 6963 3410 7010 3428
rect 6963 3383 6979 3410
rect 7000 3383 7010 3410
rect 6963 3113 7010 3383
rect 6963 3086 6974 3113
rect 6995 3086 7010 3113
rect 6963 3068 7010 3086
rect 17118 3315 17142 3334
rect 17118 3295 17121 3315
rect 17138 3295 17142 3315
rect 17118 3114 17142 3295
rect 17118 3093 17121 3114
rect 17138 3093 17142 3114
rect 17118 3085 17142 3093
rect 5401 1937 5444 1955
rect 5401 1913 5421 1937
rect 5441 1913 5444 1937
rect 5401 1769 5444 1913
rect 5401 1745 5408 1769
rect 5428 1745 5444 1769
rect 5401 1740 5444 1745
rect 15507 1925 15569 1943
rect 15507 1892 15529 1925
rect 15552 1892 15569 1925
rect 15507 1709 15569 1892
rect 15507 1676 15532 1709
rect 15555 1676 15569 1709
rect 15507 1664 15569 1676
rect 3741 1063 3775 1078
rect 3741 1035 3746 1063
rect 3764 1035 3775 1063
rect 3741 875 3775 1035
rect 3741 847 3746 875
rect 3764 847 3775 875
rect 3741 840 3775 847
rect 13883 1051 13927 1086
rect 13883 1016 13897 1051
rect 13923 1016 13927 1051
rect 13883 815 13927 1016
rect 13883 780 13888 815
rect 13914 780 13927 815
rect 13883 772 13927 780
rect 12110 626 12164 656
rect 1985 602 2020 613
rect 1985 583 1995 602
rect 2017 583 2020 602
rect 1985 507 2020 583
rect 1985 488 1993 507
rect 2015 488 2020 507
rect 1985 482 2020 488
rect 12110 596 12138 626
rect 12161 596 12164 626
rect 12110 464 12164 596
rect 12110 434 12132 464
rect 12155 434 12164 464
rect 12110 428 12164 434
rect 472 302 504 307
rect 468 299 504 302
rect 468 280 474 299
rect 496 280 504 299
rect 468 263 504 280
rect 10594 288 10631 296
rect 10594 263 10603 288
rect 10621 263 10631 288
rect 468 259 505 263
rect 466 237 510 259
rect 466 235 506 237
rect 475 212 506 235
rect 472 206 506 212
rect 472 204 509 206
rect 472 185 479 204
rect 501 185 509 204
rect 472 182 509 185
rect 10594 183 10631 263
rect 472 181 505 182
rect 10594 158 10603 183
rect 10621 158 10631 183
rect 10594 156 10631 158
rect 10594 153 10630 156
rect 13856 -440 13904 -414
rect 12118 -460 12149 -446
rect 10603 -483 10634 -476
rect 10603 -500 10608 -483
rect 10625 -500 10634 -483
rect 10603 -503 10634 -500
rect 12118 -486 12124 -460
rect 12145 -486 12149 -460
rect 13856 -469 13862 -440
rect 13888 -442 13904 -440
rect 15524 -415 15588 -401
rect 13888 -469 13906 -442
rect 13856 -481 13906 -469
rect 10604 -1195 10622 -503
rect 12118 -1138 12149 -486
rect 13857 -1020 13906 -481
rect 15524 -457 15540 -415
rect 15578 -457 15588 -415
rect 15524 -829 15588 -457
rect 17097 -449 17140 -438
rect 17097 -470 17107 -449
rect 17130 -470 17140 -449
rect 17097 -741 17140 -470
rect 17097 -762 17109 -741
rect 17132 -762 17140 -741
rect 17097 -806 17140 -762
rect 15524 -871 15586 -829
rect 15524 -913 15530 -871
rect 15568 -913 15586 -871
rect 15524 -927 15586 -913
rect 13857 -1049 13870 -1020
rect 13896 -1049 13906 -1020
rect 13857 -1059 13906 -1049
rect 12118 -1163 12125 -1138
rect 12121 -1164 12125 -1163
rect 12146 -1164 12149 -1138
rect 12121 -1173 12149 -1164
rect 10600 -1202 10630 -1195
rect 10600 -1220 10605 -1202
rect 10623 -1220 10630 -1202
rect 10600 -1226 10630 -1220
<< via1 >>
rect 21904 12662 21933 12690
rect 21530 12276 21559 12306
<< metal2 >>
rect 9569 24232 12052 24235
rect 8175 24230 12052 24232
rect 5384 24192 12052 24230
rect 5384 24189 9593 24192
rect 5384 24187 8198 24189
rect 5384 21799 5416 24187
rect 12030 24181 12052 24192
rect 12030 23881 12058 24181
rect 12030 23254 12063 23881
rect 12030 23235 12066 23254
rect 12033 22608 12066 23235
rect 5384 21759 5427 21799
rect 5389 21010 5427 21759
rect 21896 12732 21943 12741
rect 21896 12704 21904 12732
rect 21933 12704 21943 12732
rect 21896 12690 21943 12704
rect 21896 12662 21904 12690
rect 21933 12662 21943 12690
rect 21896 12658 21943 12662
rect 21475 12310 21564 12312
rect 21472 12306 21564 12310
rect 21472 12276 21530 12306
rect 21559 12276 21564 12306
rect 21472 12263 21564 12276
rect 21472 11917 21490 12263
rect 18600 11895 20985 11901
rect 21472 11895 21488 11917
rect 18600 11878 21488 11895
rect 21472 11877 21488 11878
<< via2 >>
rect 21904 12704 21933 12732
<< metal3 >>
rect 21895 12784 21945 12787
rect 21895 12750 21905 12784
rect 21938 12750 21945 12784
rect 21895 12732 21945 12750
rect 21895 12704 21904 12732
rect 21933 12704 21945 12732
rect 21895 12699 21945 12704
<< via3 >>
rect 21905 12750 21938 12784
<< metal4 >>
rect 3873 24121 3921 24123
rect 11230 24121 11295 24123
rect 3873 24080 11295 24121
rect 3873 23743 3921 24080
rect 11230 24079 11295 24080
rect 11257 23912 11295 24079
rect 19270 13119 21319 13120
rect 21894 13119 21942 13120
rect 19270 13085 21942 13119
rect 19270 13082 21319 13085
rect 21894 12813 21942 13085
rect 21894 12806 21945 12813
rect 21895 12784 21945 12806
rect 21895 12750 21905 12784
rect 21938 12750 21945 12784
rect 21895 12747 21945 12750
use 6bitdac_layout  6bitdac_layout_0
timestamp 1616477680
transform 1 0 122 0 1 12065
box -122 -12065 9858 11921
use 6bitdac_layout  6bitdac_layout_1
timestamp 1616477680
transform 1 0 10253 0 1 12046
box -122 -12065 9858 11921
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 21448 0 1 12168
box 20 86 1230 590
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 -88 0 1 -10
box 109 -171 242 -45
<< labels >>
rlabel locali 43 -58 43 -58 1 x1_vref5
rlabel locali 127 -201 127 -201 1 x2_vref1
rlabel locali 10218 -44 10218 -44 1 inp2
rlabel locali 287 23972 287 23972 1 inp1
rlabel locali 21457 12444 21457 12445 1 d6
rlabel locali 22712 12530 22712 12530 1 out_v
rlabel metal4 21921 12796 21921 12796 1 vdd!
rlabel metal2 21500 12279 21500 12279 1 gnd!
rlabel locali 22598 12148 22598 12148 1 x2_out_v
rlabel locali 22577 12816 22577 12816 1 x1_out_v
rlabel locali 489 127 489 127 1 d0
rlabel locali 1996 107 1996 107 1 d1
rlabel locali 5426 240 5426 240 1 d3
rlabel locali 7001 463 7001 463 1 d4
rlabel locali 8663 405 8663 405 1 d5
rlabel locali 3743 -587 3743 -587 1 d2
<< end >>
