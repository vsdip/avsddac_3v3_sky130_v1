magic
tech sky130A
magscale 1 2
timestamp 1624910849
<< locali >>
rect 1224 111478 1280 111678
rect 166990 55698 167030 58214
rect 170054 56858 170108 57650
rect 173560 56638 173644 58478
rect 176982 54874 177048 58546
rect 179826 56758 179890 57852
rect 183168 54830 183216 58556
rect 188400 54802 188470 58594
rect 191890 54838 191964 58672
rect 196096 54788 196172 79662
rect 205436 57549 205476 57550
rect 205436 57515 205439 57549
rect 205473 57515 205476 57549
rect 205436 57514 205476 57515
rect 202790 57336 203012 57432
rect 166000 5276 166054 5432
<< viali >>
rect 205439 57515 205473 57549
<< metal1 >>
rect 205430 57564 205602 57576
rect 205430 57549 205547 57564
rect 205430 57515 205439 57549
rect 205473 57515 205547 57549
rect 205430 57512 205547 57515
rect 205599 57512 205602 57564
rect 205430 57500 205602 57512
rect 208338 52576 208562 52648
<< via1 >>
rect 205547 57512 205599 57564
<< metal2 >>
rect 196548 55424 196626 85814
rect 205538 57568 205722 57578
rect 205538 57564 205651 57568
rect 205538 57512 205547 57564
rect 205599 57512 205651 57564
rect 205707 57512 205722 57568
rect 205538 57500 205722 57512
<< via2 >>
rect 205651 57512 205707 57568
<< metal3 >>
rect 205750 57584 205862 57590
rect 205638 57576 205862 57584
rect 205638 57568 205771 57576
rect 205638 57512 205651 57568
rect 205707 57512 205771 57568
rect 205835 57512 205862 57576
rect 205638 57500 205862 57512
rect 205750 57498 205862 57500
rect 207214 49908 236658 79834
<< via3 >>
rect 205771 57512 205835 57576
<< mimcap >>
rect 208484 57576 235206 78746
rect 208484 57512 210209 57576
rect 210273 57512 235206 57576
rect 208484 51540 235206 57512
<< mimcapcontact >>
rect 210209 57512 210273 57576
<< metal4 >>
rect 201970 58220 202162 83072
rect 205764 57576 210286 57584
rect 205764 57512 205771 57576
rect 205835 57512 210209 57576
rect 210273 57512 210286 57576
rect 205764 57504 210286 57512
rect 205764 57500 205956 57504
use cap_28p  cap_28p_0
timestamp 1624819264
transform 1 0 210498 0 1 53878
box -1968 -2452 24820 24898
use 10bitdac_layout  10bitdac_layout_0
timestamp 1624819264
transform 1 0 428 0 1 57644
box -428 -57692 205056 54770
<< labels >>
rlabel metal4 s 207420 57532 207420 57532 4 out
port 1 nsew
flabel locali s 166000 5276 166054 5432 0 FreeSans 195 0 0 0 inp2
port 2 nsew
flabel locali s 1224 111478 1280 111678 0 FreeSans 195 0 0 0 inp1
port 3 nsew
flabel locali s 166990 55698 167030 58214 0 FreeSans 195 0 0 0 d0
port 4 nsew
flabel locali s 170054 56858 170108 57650 0 FreeSans 195 0 0 0 d1
port 5 nsew
flabel locali s 173560 56638 173644 58478 0 FreeSans 195 0 0 0 d2
port 6 nsew
flabel locali s 176982 54874 177048 58546 0 FreeSans 195 0 0 0 d3
port 7 nsew
flabel locali s 179826 56758 179890 57852 0 FreeSans 195 0 0 0 d4
port 8 nsew
flabel locali s 183168 54830 183216 58556 0 FreeSans 195 0 0 0 d5
port 9 nsew
flabel locali s 188400 54802 188470 58594 0 FreeSans 195 0 0 0 d6
port 10 nsew
flabel locali s 191890 54838 191964 58672 0 FreeSans 195 0 0 0 d7
port 11 nsew
flabel locali s 196096 54788 196172 79662 0 FreeSans 195 0 0 0 d8
port 12 nsew
flabel locali s 202790 57336 203012 57432 0 FreeSans 195 0 0 0 d9
port 13 nsew
flabel metal2 s 196548 55424 196626 85814 0 FreeSans 195 0 0 0 gnd!
port 14 nsew
flabel metal4 s 201970 58220 202162 83072 0 FreeSans 195 0 0 0 vdd!
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 1748 1088
<< end >>
