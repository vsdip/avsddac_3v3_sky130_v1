magic
tech sky130A
timestamp 1616475377
<< locali >>
rect 90 1091 116 1186
rect 4390 775 4837 778
rect 3296 772 4837 775
rect 3229 737 4837 772
rect 3229 734 4427 737
rect 3229 733 3318 734
rect 1919 480 1969 707
rect 1919 462 1932 480
rect 1955 462 1969 480
rect 1919 442 1969 462
rect 4799 351 4835 737
rect 371 137 419 284
rect 371 115 383 137
rect 402 115 419 137
rect 371 99 419 115
rect 1901 262 1967 271
rect 1901 244 1932 262
rect 1955 244 1967 262
rect 0 -9 104 8
rect 85 -139 104 -9
rect -27 -306 -8 -180
rect 373 -247 419 -238
rect 373 -269 387 -247
rect 406 -269 419 -247
rect 73 -306 100 -305
rect -27 -327 100 -306
rect 73 -348 100 -327
rect 373 -312 419 -269
rect 1901 -311 1967 244
rect 4893 210 5060 217
rect 4893 190 4901 210
rect 4921 190 5060 210
rect 4893 186 5060 190
rect 3674 104 3747 150
rect 373 -497 421 -312
rect 1901 -329 1916 -311
rect 1939 -329 1967 -311
rect 1901 -342 1967 -329
rect 1904 -526 1954 -519
rect 1904 -544 1917 -526
rect 1940 -544 1954 -526
rect 1904 -784 1954 -544
rect 4820 -667 4854 -18
rect 4763 -669 4859 -667
rect 3211 -671 3639 -670
rect 4379 -671 4859 -669
rect 3211 -703 4859 -671
rect 3211 -704 4425 -703
rect 3610 -705 4425 -704
rect 4763 -707 4859 -703
rect 4820 -708 4854 -707
rect -16 -1468 10 -1409
rect -18 -1530 12 -1468
<< viali >>
rect 1932 462 1955 480
rect 383 115 402 137
rect 1932 244 1955 262
rect 387 -269 406 -247
rect 4901 190 4921 210
rect 1916 -329 1939 -311
rect 1917 -544 1940 -526
<< metal1 >>
rect 1917 480 1967 497
rect 1917 462 1932 480
rect 1955 462 1967 480
rect 1917 262 1967 462
rect 4136 370 4189 376
rect 4136 338 4149 370
rect 4182 338 4189 370
rect 4136 335 4189 338
rect 1917 244 1932 262
rect 1955 244 1967 262
rect 1917 232 1967 244
rect 371 137 420 145
rect 371 115 383 137
rect 402 115 420 137
rect 371 -247 420 115
rect 3779 -15 3817 8
rect 3779 -51 3783 -15
rect 3815 -51 3817 -15
rect 3779 -64 3817 -51
rect 371 -269 387 -247
rect 406 -269 420 -247
rect 371 -278 420 -269
rect 1902 -311 1952 -300
rect 1902 -329 1916 -311
rect 1939 -329 1952 -311
rect 1902 -526 1952 -329
rect 1902 -544 1917 -526
rect 1940 -544 1952 -526
rect 1902 -565 1952 -544
<< via1 >>
rect 4149 338 4182 370
rect 3783 -51 3815 -15
<< metal2 >>
rect 4145 414 4190 421
rect 4145 381 4151 414
rect 4182 381 4190 414
rect 4145 370 4190 381
rect 4145 338 4149 370
rect 4182 338 4190 370
rect 4145 335 4190 338
rect 1728 -641 1753 -3
rect 3714 -11 3819 -9
rect 3713 -15 3819 -11
rect 3713 -51 3783 -15
rect 3815 -51 3819 -15
rect 3713 -61 3819 -51
rect 3713 -136 3745 -61
rect 3713 -293 3744 -136
rect 1725 -1479 1755 -641
rect 3710 -1383 3746 -293
rect 2534 -1420 3411 -1419
rect 3710 -1420 3743 -1383
rect 2534 -1425 3743 -1420
rect 2448 -1426 3743 -1425
rect 2146 -1427 3743 -1426
rect 1940 -1448 3743 -1427
rect 1940 -1449 2555 -1448
rect 3381 -1449 3743 -1448
rect 1940 -1450 2456 -1449
rect 1940 -1451 2149 -1450
<< via2 >>
rect 4151 381 4182 414
<< metal3 >>
rect 4145 487 4190 494
rect 4145 454 4151 487
rect 4185 454 4190 487
rect 4145 414 4190 454
rect 4145 381 4151 414
rect 4182 381 4190 414
rect 4145 377 4190 381
<< via3 >>
rect 4151 454 4185 487
<< metal4 >>
rect 3387 1135 3438 1148
rect 3860 1135 4193 1137
rect 3170 1132 4193 1135
rect 3114 1131 4193 1132
rect 2943 1130 4193 1131
rect 2434 1095 4193 1130
rect 2434 1094 3121 1095
rect 2434 1093 2950 1094
rect 3170 1091 4193 1095
rect 3387 -57 3438 1091
rect 3860 1087 4193 1091
rect 4146 512 4190 1087
rect 4145 487 4190 512
rect 4145 454 4151 487
rect 4185 454 4190 487
rect 4145 450 4190 454
rect 3387 -88 3436 -57
rect 2719 -108 3436 -88
rect 2365 -166 3436 -108
rect 2365 -168 2747 -166
use 2bitdac_layout  2bitdac_layout_1
timestamp 1616473885
transform 1 0 -12 0 1 -825
box -5 -649 3251 715
use 2bitdac_layout  2bitdac_layout_0
timestamp 1616473885
transform 1 0 5 0 1 617
box -5 -649 3251 715
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 3697 0 1 -155
box 20 86 1230 590
use res250_layout  res250_layout_0
timestamp 1615764517
transform 0 1 148 -1 0 14
box 109 -171 242 -45
<< labels >>
rlabel locali -1 -1455 -1 -1455 1 inp2
rlabel locali 103 1153 103 1153 1 inp1
rlabel locali 92 -76 92 -76 1 x1_vref5
rlabel locali -20 -259 -20 -259 1 x2_vref1
rlabel locali 399 -353 399 -353 1 d0
rlabel locali 1919 -53 1919 -53 1 d1
rlabel locali 3706 134 3706 134 1 d2
rlabel locali 3352 755 3352 755 1 x1_out_v
rlabel locali 3292 -685 3292 -685 1 x2_out_v
rlabel locali 4993 200 4993 200 1 out_v
rlabel metal4 3773 1113 3773 1113 1 vdd!
rlabel metal2 3731 -1350 3731 -1350 1 gnd!
<< end >>
