magic
tech sky130A
magscale 1 2
timestamp 1624221218
<< checkpaint >>
rect -1314 -4320 11380 3924
<< locali >>
rect 180 2182 232 2372
rect 8780 1550 9674 1556
rect 6592 1544 9674 1550
rect 6458 1474 9674 1544
rect 6458 1468 8854 1474
rect 6458 1466 6636 1468
rect 3838 959 3938 1414
rect 3838 925 3870 959
rect 3904 925 3938 959
rect 3838 884 3938 925
rect 9598 702 9670 1474
rect 742 269 838 568
rect 742 235 768 269
rect 802 235 838 269
rect 742 198 838 235
rect 3802 523 3934 542
rect 3802 489 3870 523
rect 3904 489 3934 523
rect 0 -18 208 16
rect 170 -278 208 -18
rect -54 -612 -16 -360
rect 746 -499 838 -476
rect 746 -533 776 -499
rect 810 -533 838 -499
rect 146 -612 200 -610
rect -54 -654 200 -612
rect 146 -696 200 -654
rect 746 -624 838 -533
rect 3802 -623 3934 489
rect 9786 417 10120 434
rect 9786 383 9805 417
rect 9839 383 10120 417
rect 9786 372 10120 383
rect 7348 208 7494 300
rect 746 -994 842 -624
rect 3802 -657 3838 -623
rect 3872 -657 3934 -623
rect 3802 -684 3934 -657
rect 3808 -1053 3908 -1038
rect 3808 -1087 3840 -1053
rect 3874 -1087 3908 -1053
rect 3808 -1568 3908 -1087
rect 9640 -1334 9708 -36
rect 9526 -1338 9718 -1334
rect 6422 -1342 7278 -1340
rect 8758 -1342 9718 -1338
rect 6422 -1406 9718 -1342
rect 6422 -1408 8850 -1406
rect 7220 -1410 8850 -1408
rect 9526 -1414 9718 -1406
rect 9640 -1416 9708 -1414
rect -32 -2936 20 -2818
rect -36 -3060 24 -2936
<< viali >>
rect 3870 925 3904 959
rect 768 235 802 269
rect 3870 489 3904 523
rect 776 -533 810 -499
rect 9805 383 9839 417
rect 3838 -657 3872 -623
rect 3840 -1087 3874 -1053
<< metal1 >>
rect 3834 959 3934 994
rect 3834 925 3870 959
rect 3904 925 3934 959
rect 3834 523 3934 925
rect 8272 734 8378 752
rect 8272 682 8305 734
rect 8357 682 8378 734
rect 8272 670 8378 682
rect 3834 489 3870 523
rect 3904 489 3934 523
rect 3834 464 3934 489
rect 9802 417 9842 420
rect 9802 383 9805 417
rect 9839 383 9842 417
rect 9802 380 9842 383
rect 742 269 840 290
rect 742 235 768 269
rect 802 235 840 269
rect 742 -499 840 235
rect 7558 -40 7634 16
rect 7558 -92 7572 -40
rect 7624 -92 7634 -40
rect 7558 -128 7634 -92
rect 742 -533 776 -499
rect 810 -533 840 -499
rect 742 -556 840 -533
rect 3804 -623 3904 -600
rect 3804 -657 3838 -623
rect 3872 -657 3904 -623
rect 3804 -1053 3904 -657
rect 3804 -1087 3840 -1053
rect 3874 -1087 3904 -1053
rect 3804 -1130 3904 -1087
<< via1 >>
rect 8305 682 8357 734
rect 7572 -92 7624 -40
<< metal2 >>
rect 8290 823 8380 842
rect 8290 767 8305 823
rect 8361 767 8380 823
rect 8290 734 8380 767
rect 8290 682 8305 734
rect 8357 682 8380 734
rect 8290 670 8380 682
rect 3456 -1282 3506 -6
rect 7428 -22 7638 -18
rect 7426 -40 7638 -22
rect 7426 -92 7572 -40
rect 7624 -92 7638 -40
rect 7426 -122 7638 -92
rect 7426 -272 7490 -122
rect 7426 -586 7488 -272
rect 3450 -2958 3510 -1282
rect 7420 -2766 7492 -586
rect 5068 -2840 6822 -2838
rect 7420 -2840 7486 -2766
rect 5068 -2850 7486 -2840
rect 4896 -2852 7486 -2850
rect 4292 -2854 7486 -2852
rect 3880 -2896 7486 -2854
rect 3880 -2898 5110 -2896
rect 6762 -2898 7486 -2896
rect 3880 -2900 4912 -2898
rect 3880 -2902 4298 -2900
<< via2 >>
rect 8305 767 8361 823
<< metal3 >>
rect 8290 973 8380 988
rect 8290 909 8304 973
rect 8368 909 8380 973
rect 8290 823 8380 909
rect 8290 767 8305 823
rect 8361 767 8380 823
rect 8290 754 8380 767
<< via3 >>
rect 8304 909 8368 973
<< metal4 >>
rect 6774 2270 6876 2296
rect 7720 2270 8386 2274
rect 6340 2264 8386 2270
rect 6228 2262 8386 2264
rect 5886 2260 8386 2262
rect 4868 2190 8386 2260
rect 4868 2188 6242 2190
rect 4868 2186 5900 2188
rect 6340 2182 8386 2190
rect 6774 -114 6876 2182
rect 7720 2174 8386 2182
rect 8292 1024 8380 2174
rect 8290 973 8380 1024
rect 8290 909 8304 973
rect 8368 909 8380 973
rect 8290 900 8380 909
rect 6774 -176 6872 -114
rect 5438 -216 6872 -176
rect 4730 -332 6872 -216
rect 4730 -336 5494 -332
use res250_layout  res250_layout_0
timestamp 1624221218
transform 0 1 296 -1 0 28
box 218 -342 484 -90
use switch_layout  switch_layout_0
timestamp 1624221218
transform 1 0 7394 0 1 -310
box 40 172 2460 1180
use 2bitdac_layout  2bitdac_layout_0
timestamp 1624221218
transform 1 0 10 0 1 1234
box -10 -1298 6502 1430
use 2bitdac_layout  2bitdac_layout_1
timestamp 1624221218
transform 1 0 -24 0 1 -1650
box -10 -1298 6502 1430
<< labels >>
rlabel locali s -2 -2910 -2 -2910 4 inp2
rlabel locali s 206 2306 206 2306 4 inp1
rlabel locali s 184 -152 184 -152 4 x1_vref5
rlabel locali s -40 -518 -40 -518 4 x2_vref1
rlabel locali s 798 -706 798 -706 4 d0
rlabel locali s 3838 -106 3838 -106 4 d1
rlabel locali s 7412 268 7412 268 4 d2
rlabel locali s 6704 1510 6704 1510 4 x1_out_v
rlabel locali s 6584 -1370 6584 -1370 4 x2_out_v
rlabel locali s 9986 400 9986 400 4 out_v
rlabel metal4 s 7546 2226 7546 2226 4 vdd!
rlabel metal2 s 7462 -2700 7462 -2700 4 gnd!
<< end >>
