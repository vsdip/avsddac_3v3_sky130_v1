* SPICE3 file created from 3bitdac_layout.ext - technology: sky130A

.option scale=10000u

X0 switch_layout_0/dd switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1 switch_layout_0/dd switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2 switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X3 switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X4 x1_out_v switch_layout_0/dd out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X5 out_v switch_layout_0/dinb x1_out_v switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X6 x2_out_v switch_layout_0/dd out_v switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X7 out_v switch_layout_0/dinb x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X8 2bitdac_layout_0/switch_layout_0/dd 2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X9 2bitdac_layout_0/switch_layout_0/dd 2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X10 2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X11 2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X12 2bitdac_layout_0/x1_inp1 2bitdac_layout_0/switch_layout_0/dd 2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X13 2bitdac_layout_0/x1_vout 2bitdac_layout_0/switch_layout_0/dinb 2bitdac_layout_0/x1_inp1 2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X14 2bitdac_layout_0/x1_inp2 2bitdac_layout_0/switch_layout_0/dd 2bitdac_layout_0/x1_vout 2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X15 2bitdac_layout_0/x1_vout 2bitdac_layout_0/switch_layout_0/dinb 2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X16 2bitdac_layout_0/switch_layout_1/dd 2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X17 2bitdac_layout_0/switch_layout_1/dd 2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X18 2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X19 2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X20 2bitdac_layout_0/x2_inp1 2bitdac_layout_0/switch_layout_1/dd 2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X21 2bitdac_layout_0/x2_vout 2bitdac_layout_0/switch_layout_1/dinb 2bitdac_layout_0/x2_inp1 2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X22 x1_vref5 2bitdac_layout_0/switch_layout_1/dd 2bitdac_layout_0/x2_vout 2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X23 2bitdac_layout_0/x2_vout 2bitdac_layout_0/switch_layout_1/dinb x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X24 2bitdac_layout_0/switch_layout_2/dd 2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X25 2bitdac_layout_0/switch_layout_2/dd 2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X26 2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X27 2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X28 2bitdac_layout_0/x1_vout 2bitdac_layout_0/switch_layout_2/dd x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X29 x1_out_v 2bitdac_layout_0/switch_layout_2/dinb 2bitdac_layout_0/x1_vout 2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X30 2bitdac_layout_0/x2_vout 2bitdac_layout_0/switch_layout_2/dd x1_out_v 2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X31 x1_out_v 2bitdac_layout_0/switch_layout_2/dinb 2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X32 2bitdac_layout_0/x1_inp1 2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X33 2bitdac_layout_0/x1_inp2 2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X34 inp1 2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X35 2bitdac_layout_0/x2_inp1 x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X36 2bitdac_layout_1/switch_layout_0/dd 2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X37 2bitdac_layout_1/switch_layout_0/dd 2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X38 2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X39 2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X40 2bitdac_layout_1/x1_inp1 2bitdac_layout_1/switch_layout_0/dd 2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X41 2bitdac_layout_1/x1_vout 2bitdac_layout_1/switch_layout_0/dinb 2bitdac_layout_1/x1_inp1 2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X42 2bitdac_layout_1/x1_inp2 2bitdac_layout_1/switch_layout_0/dd 2bitdac_layout_1/x1_vout 2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X43 2bitdac_layout_1/x1_vout 2bitdac_layout_1/switch_layout_0/dinb 2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X44 2bitdac_layout_1/switch_layout_1/dd 2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X45 2bitdac_layout_1/switch_layout_1/dd 2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X46 2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X47 2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X48 2bitdac_layout_1/x2_inp1 2bitdac_layout_1/switch_layout_1/dd 2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X49 2bitdac_layout_1/x2_vout 2bitdac_layout_1/switch_layout_1/dinb 2bitdac_layout_1/x2_inp1 2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X50 inp2 2bitdac_layout_1/switch_layout_1/dd 2bitdac_layout_1/x2_vout 2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X51 2bitdac_layout_1/x2_vout 2bitdac_layout_1/switch_layout_1/dinb inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X52 2bitdac_layout_1/switch_layout_2/dd 2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X53 2bitdac_layout_1/switch_layout_2/dd 2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X54 2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X55 2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X56 2bitdac_layout_1/x1_vout 2bitdac_layout_1/switch_layout_2/dd x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X57 x2_out_v 2bitdac_layout_1/switch_layout_2/dinb 2bitdac_layout_1/x1_vout 2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X58 2bitdac_layout_1/x2_vout 2bitdac_layout_1/switch_layout_2/dd x2_out_v 2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X59 x2_out_v 2bitdac_layout_1/switch_layout_2/dinb 2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X60 2bitdac_layout_1/x1_inp1 2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X61 2bitdac_layout_1/x1_inp2 2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X62 x2_vref1 2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X63 2bitdac_layout_1/x2_inp1 inp2 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X64 x1_vref5 x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
C0 vdd gnd 15.39fF
C1 d0 gnd 5.11fF
