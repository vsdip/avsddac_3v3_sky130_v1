* SPICE3 file created from 10bitdac_cap_layout_design.ext - technology: sky130A

*Model Description
.para temp =27 
.lib "../sky130_fd_pr/models/sky130.lib.spice" tt

X0 out_v 0 sky130_fd_pr__cap_mim_m3_1 l=121.48 w=120.63
X1 10bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2 10bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3 10bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d9 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4 10bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d9 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5 10bitdac_layout_0/x1_out_v 10bitdac_layout_0/switch_layout_0/dd out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6 out_v 10bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/x1_out_v 10bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7 10bitdac_layout_0/x2_out_v 10bitdac_layout_0/switch_layout_0/dd out_v 10bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8 out_v 10bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9 10bitdac_layout_0/x1_vref5 10bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X10 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X11 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X12 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d8 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X13 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X14 10bitdac_layout_0/9bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X15 10bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X16 10bitdac_layout_0/9bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X17 10bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X18 10bitdac_layout_0/9bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X19 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X20 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X21 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d7 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X22 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X23 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X24 10bitdac_layout_0/9bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X25 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X26 10bitdac_layout_0/9bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X27 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X28 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X29 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X30 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X31 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X32 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X33 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X34 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X35 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X36 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X37 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X38 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X39 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X40 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X41 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X42 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X43 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X44 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X45 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X46 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X47 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X48 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X49 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X50 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X51 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X52 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X53 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X54 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X55 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X56 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X57 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X58 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X59 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X60 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X61 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X62 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X63 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X64 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X65 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X66 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X67 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X68 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X69 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X70 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X71 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X72 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X73 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X74 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X75 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X76 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X77 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X78 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X79 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X80 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X81 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X82 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X83 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X84 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X85 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X86 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X87 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X88 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X89 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X90 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X91 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X92 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X93 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X94 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X95 10bitdac_layout_0/inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X96 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X97 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X98 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X99 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X100 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X101 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X102 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X103 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X104 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X105 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X106 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X107 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X108 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X109 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X110 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X111 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X112 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X113 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X114 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X115 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X116 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X117 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X118 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X119 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X120 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X121 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X122 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X123 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X124 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X125 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X126 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X127 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X128 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X129 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X130 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X131 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X132 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X133 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X134 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X135 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X136 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X137 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X138 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X139 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X140 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X141 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X142 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X143 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X144 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X145 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X146 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X147 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X148 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X149 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X150 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X151 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X152 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X153 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X154 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X155 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X156 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X157 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X158 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X159 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X160 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X161 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X162 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X163 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X164 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X165 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X166 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X167 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X168 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X169 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X170 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X171 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X172 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X173 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X174 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X175 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X176 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X177 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X178 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X179 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X180 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X181 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X182 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X183 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X184 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X185 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X186 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X187 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X188 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X189 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X190 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X191 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X192 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X193 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X194 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X195 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X196 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X197 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X198 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X199 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X200 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X201 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X202 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X203 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X204 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X205 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X206 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X207 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X208 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X209 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X210 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X211 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X212 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X213 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X214 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X215 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X216 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X217 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X218 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X219 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X220 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X221 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X222 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X223 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X224 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X225 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X226 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X227 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X228 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X229 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X230 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X231 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X232 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X233 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X234 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X235 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X236 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X237 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X238 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X239 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X240 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X241 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X242 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X243 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X244 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X245 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X246 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X247 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X248 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X249 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X250 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X251 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X252 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X253 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X254 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X255 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X256 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X257 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X258 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X259 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X260 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X261 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X262 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X263 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X264 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X265 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X266 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X267 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X268 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X269 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X270 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X271 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X272 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X273 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X274 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X275 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X276 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X277 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X278 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X279 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X280 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X281 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X282 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X283 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X284 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X285 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X286 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X287 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X288 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X289 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X290 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X291 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X292 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X293 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X294 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X295 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X296 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X297 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X298 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X299 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X300 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X301 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X302 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X303 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X304 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X305 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X306 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X307 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X308 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X309 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X310 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X311 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X312 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X313 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X314 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X315 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X316 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X317 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X318 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X319 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X320 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X321 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X322 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X323 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X324 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X325 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X326 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X327 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X328 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X329 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X330 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X331 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X332 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X333 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X334 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X335 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X336 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X337 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X338 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X339 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X340 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X341 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X342 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X343 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X344 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X345 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X346 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X347 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X348 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X349 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X350 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X351 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X352 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X353 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X354 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X355 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X356 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X357 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X358 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X359 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X360 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X361 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X362 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X363 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X364 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X365 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X366 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X367 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X368 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X369 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X370 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X371 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X372 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X373 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X374 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X375 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X376 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X377 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X378 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X379 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X380 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X381 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X382 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X383 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X384 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X385 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X386 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X387 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X388 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X389 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X390 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X391 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X392 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X393 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X394 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X395 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X396 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X397 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X398 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X399 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X400 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X401 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X402 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X403 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X404 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X405 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X406 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X407 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X408 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X409 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X410 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X411 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X412 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X413 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X414 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X415 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X416 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X417 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X418 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X419 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X420 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X421 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X422 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X423 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X424 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X425 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X426 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X427 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X428 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X429 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X430 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X431 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X432 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X433 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X434 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X435 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X436 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X437 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X438 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X439 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X440 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X441 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X442 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X443 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X444 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X445 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X446 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X447 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X448 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X449 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X450 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X451 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X452 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X453 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X454 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X455 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X456 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X457 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X458 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X459 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X460 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X461 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X462 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X463 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X464 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X465 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X466 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X467 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X468 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X469 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X470 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X471 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X472 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X473 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X474 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X475 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X476 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X477 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X478 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X479 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X480 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X481 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X482 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X483 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X484 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X485 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X486 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X487 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X488 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X489 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X490 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X491 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X492 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X493 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X494 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X495 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X496 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X497 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X498 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X499 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X500 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X501 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X502 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X503 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X504 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X505 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X506 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X507 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X508 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X509 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X510 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X511 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X512 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X513 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X514 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X515 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X516 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X517 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X518 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X519 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X520 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X521 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X522 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X523 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X524 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X525 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X526 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X527 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X528 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X529 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X530 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X531 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X532 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X533 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X534 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X535 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X536 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X537 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X538 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X539 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X540 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X541 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X542 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X543 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X544 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X545 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X546 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X547 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X548 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X549 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X550 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X551 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X552 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X553 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X554 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X555 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X556 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X557 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X558 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X559 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X560 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X561 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X562 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X563 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X564 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X565 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X566 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X567 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X568 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X569 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X570 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X571 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X572 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X573 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X574 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X575 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X576 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X577 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X578 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X579 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X580 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X581 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X582 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X583 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X584 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X585 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X586 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X587 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X588 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X589 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X590 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X591 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X592 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X593 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X594 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X595 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X596 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X597 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X598 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X599 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X600 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X601 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X602 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X603 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X604 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X605 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X606 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X607 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X608 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X609 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X610 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X611 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X612 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X613 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X614 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X615 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X616 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X617 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X618 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X619 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X620 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X621 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X622 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X623 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X624 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X625 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X626 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X627 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X628 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X629 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X630 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X631 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X632 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X633 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X634 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X635 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X636 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X637 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X638 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X639 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X640 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X641 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X642 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X643 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X644 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X645 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X646 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X647 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X648 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X649 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X650 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X651 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X652 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X653 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X654 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X655 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X656 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X657 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X658 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X659 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X660 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X661 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X662 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X663 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X664 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X665 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X666 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X667 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X668 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X669 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X670 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X671 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X672 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X673 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X674 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X675 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X676 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X677 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X678 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X679 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X680 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X681 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X682 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X683 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X684 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X685 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X686 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X687 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X688 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X689 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X690 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X691 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X692 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X693 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X694 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X695 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X696 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X697 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X698 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X699 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X700 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X701 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X702 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X703 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X704 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X705 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X706 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X707 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X708 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X709 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X710 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X711 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X712 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X713 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X714 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X715 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X716 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X717 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X718 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X719 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X720 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X721 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X722 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X723 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X724 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X725 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X726 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X727 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X728 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X729 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X730 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X731 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X732 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X733 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X734 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X735 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X736 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X737 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X738 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X739 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X740 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X741 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X742 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X743 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X744 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X745 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X746 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X747 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X748 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X749 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X750 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X751 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X752 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X753 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X754 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X755 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X756 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X757 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X758 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X759 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X760 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X761 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X762 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X763 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X764 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X765 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X766 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X767 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X768 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X769 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X770 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X771 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X772 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X773 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X774 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X775 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X776 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X777 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X778 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X779 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X780 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X781 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X782 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X783 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X784 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X785 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X786 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X787 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X788 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X789 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X790 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X791 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X792 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X793 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X794 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X795 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X796 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X797 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X798 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X799 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X800 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X801 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X802 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X803 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X804 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X805 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X806 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X807 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X808 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X809 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X810 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X811 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X812 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X813 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X814 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X815 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X816 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X817 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X818 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X819 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X820 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X821 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X822 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X823 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X824 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X825 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X826 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X827 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X828 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X829 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X830 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X831 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X832 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X833 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X834 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X835 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X836 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X837 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X838 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X839 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X840 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X841 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X842 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X843 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X844 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X845 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X846 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X847 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X848 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X849 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X850 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X851 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X852 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X853 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X854 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X855 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X856 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X857 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X858 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X859 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X860 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X861 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X862 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X863 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X864 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X865 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X866 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X867 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X868 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X869 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X870 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X871 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X872 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X873 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X874 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X875 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X876 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X877 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X878 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X879 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X880 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X881 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X882 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X883 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X884 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X885 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X886 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X887 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X888 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X889 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X890 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X891 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X892 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X893 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X894 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X895 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X896 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X897 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X898 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X899 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X900 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X901 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X902 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X903 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X904 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X905 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X906 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X907 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X908 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X909 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X910 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X911 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X912 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X913 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X914 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X915 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X916 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X917 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X918 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X919 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X920 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X921 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X922 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X923 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X924 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X925 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X926 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X927 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X928 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X929 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X930 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X931 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X932 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X933 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X934 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X935 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X936 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X937 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X938 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X939 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X940 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X941 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X942 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X943 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X944 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X945 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X946 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X947 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X948 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X949 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X950 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X951 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X952 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X953 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X954 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X955 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X956 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X957 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X958 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X959 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X960 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X961 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X962 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X963 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X964 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X965 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X966 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X967 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X968 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X969 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X970 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X971 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X972 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X973 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X974 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X975 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X976 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X977 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X978 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X979 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X980 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X981 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X982 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X983 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X984 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X985 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X986 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X987 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X988 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X989 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X990 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X991 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X992 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X993 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X994 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X995 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X996 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X997 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X998 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X999 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1000 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1001 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1002 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1003 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1004 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1005 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1006 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1007 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1008 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1009 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1010 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1011 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1012 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1013 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1014 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1015 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1016 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1017 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1018 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1019 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1020 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1021 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1022 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1023 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1024 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1025 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1026 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1027 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1028 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1029 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1030 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1031 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1032 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1033 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1034 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1035 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1036 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1037 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1038 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1039 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1040 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1041 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1042 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1043 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1044 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1045 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1046 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1047 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1048 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1049 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1050 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1051 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1052 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1053 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1054 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1055 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1056 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1057 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1058 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1059 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1060 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1061 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1062 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1063 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1064 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1065 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1066 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1067 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1068 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1069 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1070 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1071 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1072 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1073 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1074 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1075 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1076 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1077 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1078 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1079 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1080 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1081 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1082 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1083 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1084 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1085 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1086 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1087 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1088 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1089 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1090 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1091 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1092 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1093 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1094 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1095 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1096 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1097 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1098 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1099 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1100 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1101 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1102 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1103 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1104 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1105 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1106 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1107 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1108 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1109 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1110 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1111 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1112 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1113 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1114 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1115 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1116 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1117 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1118 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1119 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1120 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1121 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1122 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1123 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1124 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1125 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1126 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1127 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1128 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1129 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1130 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1131 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1132 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1133 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1134 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1135 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1136 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1137 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1138 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1139 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1140 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1141 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1142 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1143 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1144 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1145 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1146 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1147 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1148 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1149 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1150 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1151 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1152 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1153 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1154 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1155 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1156 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1157 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1158 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1159 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1160 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1161 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1162 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1163 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1164 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1165 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1166 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1167 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1168 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1169 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1170 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1171 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1172 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1173 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1174 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1175 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1176 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1177 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1178 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1179 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1180 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1181 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1182 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1183 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1184 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1185 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1186 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1187 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1188 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1189 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1190 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1191 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1192 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1193 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1194 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1195 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1196 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1197 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1198 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1199 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1200 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1201 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1202 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1203 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1204 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1205 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1206 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1207 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1208 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1209 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1210 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1211 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1212 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1213 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1214 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1215 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1216 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1217 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1218 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1219 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1220 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1221 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1222 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1223 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1224 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1225 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1226 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1227 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1228 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1229 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1230 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1231 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1232 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1233 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1234 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1235 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1236 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1237 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1238 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1239 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1240 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1241 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1242 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1243 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1244 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1245 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1246 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1247 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1248 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1249 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1250 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1251 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1252 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1253 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1254 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1255 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1256 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1257 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1258 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1259 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1260 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1261 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1262 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1263 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1264 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1265 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1266 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1267 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1268 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1269 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1270 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1271 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1272 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1273 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1274 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1275 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1276 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1277 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1278 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1279 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1280 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1281 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1282 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1283 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1284 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1285 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1286 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1287 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1288 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1289 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1290 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1291 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1292 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1293 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1294 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1295 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1296 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1297 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1298 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1299 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1300 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1301 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1302 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1303 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1304 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1305 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1306 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1307 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1308 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1309 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1310 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1311 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1312 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1313 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1314 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1315 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1316 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1317 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1318 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1319 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1320 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1321 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1322 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1323 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1324 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1325 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1326 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1327 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1328 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1329 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1330 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1331 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1332 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1333 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1334 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1335 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1336 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1337 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1338 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1339 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1340 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1341 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1342 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1343 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1344 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1345 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1346 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1347 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1348 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1349 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1350 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1351 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1352 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1353 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1354 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1355 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1356 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1357 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1358 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1359 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1360 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1361 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1362 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1363 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1364 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1365 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1366 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1367 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1368 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1369 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1370 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1371 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1372 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1373 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1374 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1375 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1376 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1377 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1378 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1379 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1380 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1381 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1382 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1383 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1384 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1385 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1386 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1387 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1388 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1389 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1390 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1391 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1392 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1393 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1394 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1395 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1396 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1397 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1398 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1399 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1400 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1401 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1402 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1403 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1404 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1405 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1406 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1407 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1408 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1409 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1410 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1411 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1412 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1413 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1414 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1415 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1416 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1417 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1418 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1419 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1420 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1421 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1422 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1423 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1424 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1425 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1426 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1427 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1428 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1429 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1430 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1431 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1432 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1433 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1434 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1435 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1436 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1437 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1438 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1439 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1440 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1441 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1442 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1443 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1444 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1445 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1446 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1447 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1448 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1449 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1450 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1451 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1452 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1453 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1454 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1455 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1456 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1457 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1458 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1459 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1460 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1461 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1462 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1463 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1464 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1465 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1466 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1467 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1468 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1469 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1470 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1471 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1472 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1473 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1474 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1475 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1476 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1477 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1478 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1479 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1480 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1481 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1482 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1483 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1484 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1485 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1486 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1487 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1488 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1489 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1490 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1491 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1492 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1493 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1494 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1495 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1496 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1497 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1498 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1499 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1500 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1501 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1502 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1503 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1504 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1505 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1506 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1507 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1508 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1509 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1510 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1511 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1512 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1513 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1514 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1515 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1516 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1517 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1518 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1519 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1520 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1521 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1522 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1523 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1524 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1525 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1526 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1527 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1528 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1529 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1530 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1531 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1532 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1533 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1534 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1535 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1536 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1537 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1538 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1539 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1540 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1541 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1542 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1543 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1544 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1545 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1546 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1547 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1548 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1549 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1550 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1551 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1552 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1553 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1554 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1555 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1556 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1557 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1558 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1559 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1560 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1561 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1562 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1563 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1564 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1565 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1566 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1567 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1568 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1569 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1570 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1571 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1572 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1573 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1574 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1575 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1576 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1577 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1578 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1579 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1580 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1581 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1582 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1583 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1584 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1585 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1586 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1587 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1588 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1589 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1590 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1591 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1592 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1593 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1594 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1595 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1596 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1597 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1598 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1599 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1600 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1601 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1602 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1603 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1604 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1605 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1606 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1607 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1608 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1609 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1610 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1611 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1612 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1613 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1614 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1615 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1616 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1617 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1618 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1619 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1620 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1621 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1622 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1623 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1624 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1625 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1626 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1627 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1628 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1629 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1630 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1631 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1632 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1633 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1634 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1635 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1636 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1637 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1638 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1639 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1640 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1641 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1642 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1643 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1644 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1645 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1646 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1647 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1648 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1649 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1650 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1651 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1652 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1653 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1654 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1655 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1656 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1657 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1658 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1659 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1660 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1661 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1662 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1663 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1664 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1665 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1666 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1667 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1668 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1669 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1670 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1671 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1672 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1673 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1674 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1675 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1676 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1677 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1678 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1679 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1680 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1681 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1682 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1683 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1684 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1685 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1686 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1687 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1688 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1689 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1690 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1691 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1692 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1693 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1694 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1695 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1696 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1697 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1698 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1699 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1700 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1701 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1702 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1703 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1704 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1705 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1706 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1707 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1708 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1709 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1710 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1711 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1712 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1713 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1714 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1715 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1716 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1717 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1718 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1719 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1720 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1721 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1722 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1723 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1724 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1725 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1726 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1727 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1728 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1729 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1730 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1731 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1732 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1733 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1734 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1735 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1736 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1737 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1738 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1739 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1740 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1741 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1742 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1743 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1744 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1745 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1746 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1747 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1748 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1749 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1750 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1751 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1752 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1753 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1754 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1755 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1756 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1757 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1758 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1759 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1760 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1761 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1762 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1763 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1764 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1765 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1766 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1767 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1768 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1769 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1770 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1771 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1772 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1773 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1774 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1775 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1776 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1777 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1778 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1779 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1780 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1781 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1782 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1783 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1784 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1785 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1786 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1787 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1788 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1789 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1790 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1791 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1792 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1793 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1794 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1795 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1796 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1797 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1798 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1799 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1800 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1801 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1802 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1803 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1804 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1805 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1806 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1807 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1808 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1809 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1810 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1811 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1812 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1813 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1814 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1815 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1816 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1817 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1818 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1819 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1820 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1821 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1822 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1823 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1824 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1825 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1826 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1827 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1828 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1829 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1830 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1831 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1832 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1833 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1834 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1835 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1836 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1837 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1838 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1839 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1840 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1841 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1842 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1843 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1844 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1845 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1846 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1847 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1848 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1849 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1850 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1851 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1852 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1853 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1854 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1855 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1856 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1857 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1858 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1859 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1860 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1861 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1862 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1863 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1864 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1865 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1866 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1867 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1868 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1869 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1870 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1871 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1872 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1873 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1874 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1875 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1876 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1877 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1878 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1879 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1880 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1881 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1882 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1883 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1884 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1885 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1886 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1887 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1888 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1889 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1890 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1891 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1892 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1893 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1894 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1895 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1896 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1897 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1898 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1899 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1900 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1901 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1902 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1903 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1904 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1905 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1906 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1907 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1908 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1909 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1910 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1911 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1912 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1913 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1914 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1915 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1916 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1917 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1918 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1919 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1920 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1921 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1922 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1923 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1924 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1925 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1926 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1927 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1928 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1929 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1930 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1931 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1932 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1933 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1934 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1935 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1936 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1937 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1938 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1939 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1940 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1941 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1942 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1943 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1944 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1945 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1946 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1947 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1948 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1949 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1950 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1951 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1952 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1953 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1954 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1955 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1956 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1957 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1958 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1959 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1960 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1961 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1962 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1963 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1964 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1965 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1966 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1967 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1968 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1969 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1970 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1971 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1972 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1973 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1974 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1975 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1976 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1977 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1978 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1979 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1980 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1981 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1982 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1983 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1984 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1985 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1986 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1987 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1988 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1989 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1990 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1991 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1992 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1993 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1994 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1995 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1996 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1997 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1998 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1999 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2000 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2001 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2002 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2003 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2004 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2005 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2006 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2007 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2008 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2009 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2010 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2011 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2012 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2013 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2014 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2015 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2016 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2017 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2018 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2019 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2020 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2021 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2022 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2023 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2024 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2025 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2026 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2027 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2028 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2029 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2030 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2031 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2032 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2033 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2034 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2035 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2036 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2037 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2038 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2039 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2040 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2041 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2042 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2043 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2044 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2045 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2046 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2047 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2048 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2049 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2050 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2051 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2052 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2053 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2054 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2055 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2056 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2057 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2058 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2059 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2060 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2061 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2062 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2063 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2064 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2065 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2066 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2067 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2068 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2069 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2070 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2071 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2072 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2073 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2074 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2075 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2076 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2077 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2078 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2079 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2080 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2081 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2082 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2083 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2084 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2085 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2086 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2087 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2088 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2089 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2090 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2091 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2092 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2093 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2094 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2095 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2096 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2097 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2098 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2099 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2100 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2101 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2102 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2103 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2104 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2105 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2106 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2107 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2108 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2109 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2110 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2111 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2112 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2113 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2114 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2115 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2116 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2117 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2118 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2119 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2120 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2121 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2122 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2123 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2124 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2125 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2126 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2127 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2128 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2129 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2130 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2131 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2132 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2133 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2134 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2135 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2136 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2137 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2138 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2139 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2140 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2141 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2142 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2143 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2144 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2145 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2146 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2147 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2148 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2149 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2150 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2151 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2152 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2153 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2154 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2155 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2156 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2157 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2158 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2159 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2160 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2161 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2162 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2163 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2164 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2165 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2166 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2167 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2168 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2169 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2170 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2171 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2172 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2173 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2174 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2175 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2176 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2177 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2178 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2179 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2180 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2181 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2182 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2183 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2184 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2185 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2186 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2187 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2188 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2189 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2190 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2191 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2192 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2193 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2194 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2195 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2196 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2197 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2198 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2199 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2200 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2201 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2202 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2203 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2204 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2205 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2206 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2207 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2208 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2209 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2210 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2211 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2212 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2213 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2214 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2215 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2216 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2217 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2218 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2219 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2220 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2221 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2222 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2223 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2224 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2225 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2226 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2227 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2228 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2229 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2230 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2231 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2232 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2233 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2234 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2235 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2236 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2237 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2238 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2239 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2240 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2241 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2242 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2243 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2244 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2245 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2246 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2247 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2248 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2249 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2250 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2251 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2252 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2253 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2254 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2255 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2256 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2257 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2258 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2259 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2260 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2261 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2262 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2263 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2264 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2265 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2266 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2267 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2268 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2269 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2270 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2271 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2272 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2273 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2274 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2275 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2276 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2277 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2278 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2279 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2280 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2281 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2282 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2283 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2284 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2285 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2286 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2287 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2288 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2289 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2290 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2291 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2292 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2293 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2294 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2295 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2296 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2297 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2298 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2299 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2300 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2301 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2302 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2303 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2304 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2305 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2306 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2307 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2308 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2309 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2310 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2311 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2312 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2313 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2314 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2315 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2316 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2317 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2318 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2319 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2320 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2321 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2322 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2323 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2324 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2325 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2326 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2327 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2328 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2329 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2330 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2331 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2332 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2333 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2334 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2335 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2336 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2337 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2338 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2339 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2340 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2341 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2342 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2343 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2344 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2345 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2346 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2347 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2348 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2349 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2350 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2351 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2352 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2353 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2354 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2355 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2356 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2357 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2358 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2359 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2360 10bitdac_layout_0/9bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2361 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2362 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2363 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2364 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2365 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2366 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2367 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2368 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2369 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2370 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2371 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2372 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2373 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2374 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2375 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2376 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2377 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2378 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2379 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2380 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d7 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2381 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2382 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2383 10bitdac_layout_0/9bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2384 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2385 10bitdac_layout_0/9bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2386 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2387 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2388 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2389 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2390 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2391 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2392 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2393 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2394 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2395 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2396 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2397 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2398 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2399 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2400 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2401 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2402 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2403 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2404 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2405 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2406 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2407 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2408 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2409 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2410 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2411 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2412 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2413 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2414 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2415 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2416 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2417 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2418 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2419 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2420 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2421 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2422 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2423 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2424 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2425 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2426 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2427 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2428 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2429 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2430 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2431 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2432 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2433 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2434 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2435 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2436 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2437 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2438 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2439 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2440 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2441 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2442 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2443 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2444 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2445 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2446 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2447 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2448 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2449 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2450 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2451 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2452 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2453 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2454 10bitdac_layout_0/9bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2455 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2456 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2457 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2458 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2459 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2460 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2461 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2462 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2463 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2464 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2465 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2466 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2467 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2468 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2469 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2470 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2471 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2472 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2473 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2474 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2475 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2476 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2477 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2478 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2479 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2480 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2481 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2482 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2483 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2484 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2485 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2486 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2487 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2488 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2489 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2490 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2491 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2492 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2493 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2494 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2495 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2496 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2497 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2498 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2499 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2500 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2501 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2502 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2503 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2504 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2505 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2506 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2507 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2508 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2509 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2510 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2511 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2512 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2513 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2514 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2515 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2516 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2517 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2518 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2519 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2520 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2521 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2522 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2523 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2524 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2525 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2526 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2527 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2528 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2529 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2530 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2531 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2532 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2533 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2534 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2535 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2536 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2537 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2538 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2539 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2540 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2541 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2542 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2543 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2544 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2545 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2546 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2547 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2548 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2549 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2550 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2551 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2552 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2553 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2554 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2555 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2556 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2557 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2558 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2559 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2560 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2561 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2562 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2563 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2564 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2565 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2566 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2567 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2568 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2569 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2570 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2571 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2572 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2573 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2574 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2575 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2576 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2577 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2578 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2579 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2580 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2581 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2582 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2583 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2584 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2585 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2586 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2587 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2588 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2589 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2590 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2591 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2592 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2593 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2594 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2595 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2596 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2597 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2598 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2599 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2600 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2601 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2602 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2603 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2604 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2605 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2606 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2607 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2608 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2609 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2610 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2611 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2612 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2613 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2614 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2615 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2616 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2617 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2618 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2619 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2620 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2621 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2622 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2623 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2624 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2625 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2626 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2627 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2628 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2629 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2630 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2631 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2632 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2633 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2634 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2635 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2636 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2637 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2638 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2639 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2640 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2641 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2642 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2643 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2644 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2645 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2646 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2647 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2648 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2649 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2650 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2651 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2652 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2653 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2654 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2655 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2656 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2657 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2658 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2659 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2660 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2661 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2662 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2663 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2664 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2665 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2666 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2667 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2668 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2669 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2670 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2671 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2672 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2673 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2674 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2675 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2676 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2677 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2678 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2679 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2680 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2681 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2682 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2683 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2684 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2685 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2686 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2687 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2688 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2689 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2690 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2691 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2692 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2693 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2694 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2695 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2696 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2697 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2698 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2699 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2700 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2701 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2702 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2703 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2704 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2705 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2706 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2707 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2708 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2709 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2710 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2711 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2712 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2713 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2714 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2715 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2716 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2717 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2718 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2719 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2720 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2721 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2722 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2723 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2724 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2725 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2726 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2727 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2728 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2729 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2730 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2731 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2732 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2733 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2734 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2735 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2736 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2737 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2738 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2739 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2740 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2741 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2742 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2743 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2744 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2745 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2746 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2747 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2748 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2749 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2750 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2751 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2752 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2753 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2754 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2755 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2756 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2757 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2758 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2759 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2760 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2761 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2762 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2763 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2764 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2765 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2766 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2767 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2768 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2769 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2770 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2771 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2772 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2773 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2774 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2775 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2776 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2777 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2778 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2779 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2780 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2781 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2782 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2783 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2784 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2785 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2786 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2787 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2788 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2789 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2790 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2791 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2792 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2793 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2794 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2795 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2796 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2797 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2798 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2799 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2800 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2801 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2802 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2803 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2804 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2805 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2806 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2807 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2808 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2809 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2810 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2811 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2812 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2813 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2814 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2815 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2816 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2817 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2818 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2819 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2820 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2821 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2822 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2823 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2824 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2825 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2826 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2827 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2828 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2829 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2830 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2831 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2832 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2833 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2834 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2835 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2836 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2837 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2838 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2839 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2840 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2841 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2842 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2843 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2844 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2845 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2846 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2847 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2848 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2849 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2850 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2851 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2852 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2853 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2854 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2855 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2856 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2857 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2858 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2859 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2860 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2861 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2862 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2863 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2864 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2865 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2866 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2867 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2868 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2869 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2870 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2871 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2872 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2873 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2874 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2875 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2876 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2877 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2878 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2879 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2880 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2881 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2882 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2883 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2884 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2885 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2886 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2887 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2888 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2889 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2890 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2891 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2892 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2893 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2894 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2895 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2896 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2897 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2898 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2899 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2900 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2901 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2902 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2903 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2904 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2905 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2906 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2907 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2908 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2909 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2910 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2911 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2912 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2913 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2914 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2915 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2916 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2917 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2918 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2919 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2920 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2921 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2922 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2923 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2924 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2925 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2926 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2927 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2928 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2929 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2930 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2931 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2932 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2933 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2934 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2935 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2936 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2937 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2938 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2939 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2940 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2941 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2942 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2943 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2944 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2945 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2946 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2947 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2948 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2949 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2950 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2951 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2952 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2953 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2954 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2955 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2956 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2957 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2958 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2959 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2960 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2961 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2962 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2963 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2964 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2965 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2966 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2967 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2968 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2969 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2970 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2971 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2972 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2973 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2974 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2975 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2976 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2977 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2978 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2979 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2980 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2981 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2982 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2983 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2984 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2985 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2986 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2987 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2988 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2989 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2990 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2991 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2992 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2993 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2994 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2995 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2996 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2997 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2998 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2999 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3000 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3001 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3002 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3003 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3004 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3005 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3006 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3007 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3008 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3009 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3010 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3011 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3012 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3013 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3014 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3015 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3016 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3017 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3018 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3019 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3020 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3021 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3022 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3023 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3024 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3025 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3026 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3027 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3028 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3029 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3030 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3031 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3032 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3033 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3034 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3035 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3036 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3037 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3038 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3039 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3040 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3041 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3042 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3043 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3044 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3045 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3046 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3047 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3048 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3049 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3050 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3051 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3052 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3053 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3054 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3055 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3056 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3057 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3058 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3059 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3060 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3061 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3062 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3063 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3064 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3065 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3066 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3067 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3068 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3069 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3070 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3071 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3072 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3073 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3074 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3075 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3076 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3077 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3078 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3079 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3080 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3081 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3082 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3083 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3084 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3085 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3086 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3087 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3088 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3089 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3090 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3091 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3092 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3093 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3094 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3095 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3096 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3097 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3098 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3099 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3100 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3101 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3102 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3103 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3104 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3105 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3106 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3107 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3108 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3109 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3110 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3111 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3112 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3113 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3114 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3115 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3116 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3117 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3118 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3119 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3120 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3121 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3122 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3123 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3124 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3125 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3126 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3127 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3128 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3129 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3130 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3131 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3132 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3133 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3134 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3135 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3136 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3137 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3138 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3139 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3140 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3141 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3142 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3143 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3144 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3145 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3146 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3147 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3148 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3149 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3150 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3151 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3152 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3153 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3154 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3155 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3156 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3157 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3158 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3159 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3160 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3161 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3162 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3163 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3164 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3165 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3166 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3167 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3168 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3169 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3170 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3171 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3172 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3173 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3174 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3175 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3176 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3177 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3178 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3179 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3180 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3181 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3182 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3183 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3184 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3185 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3186 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3187 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3188 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3189 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3190 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3191 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3192 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3193 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3194 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3195 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3196 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3197 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3198 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3199 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3200 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3201 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3202 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3203 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3204 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3205 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3206 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3207 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3208 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3209 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3210 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3211 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3212 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3213 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3214 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3215 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3216 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3217 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3218 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3219 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3220 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3221 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3222 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3223 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3224 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3225 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3226 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3227 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3228 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3229 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3230 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3231 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3232 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3233 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3234 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3235 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3236 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3237 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3238 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3239 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3240 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3241 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3242 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3243 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3244 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3245 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3246 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3247 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3248 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3249 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3250 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3251 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3252 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3253 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3254 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3255 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3256 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3257 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3258 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3259 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3260 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3261 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3262 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3263 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3264 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3265 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3266 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3267 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3268 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3269 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3270 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3271 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3272 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3273 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3274 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3275 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3276 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3277 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3278 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3279 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3280 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3281 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3282 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3283 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3284 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3285 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3286 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3287 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3288 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3289 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3290 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3291 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3292 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3293 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3294 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3295 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3296 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3297 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3298 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3299 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3300 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3301 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3302 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3303 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3304 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3305 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3306 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3307 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3308 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3309 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3310 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3311 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3312 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3313 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3314 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3315 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3316 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3317 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3318 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3319 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3320 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3321 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3322 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3323 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3324 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3325 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3326 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3327 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3328 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3329 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3330 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3331 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3332 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3333 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3334 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3335 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3336 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3337 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3338 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3339 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3340 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3341 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3342 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3343 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3344 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3345 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3346 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3347 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3348 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3349 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3350 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3351 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3352 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3353 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3354 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3355 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3356 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3357 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3358 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3359 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3360 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3361 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3362 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3363 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3364 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3365 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3366 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3367 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3368 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3369 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3370 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3371 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3372 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3373 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3374 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3375 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3376 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3377 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3378 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3379 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3380 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3381 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3382 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3383 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3384 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3385 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3386 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3387 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3388 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3389 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3390 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3391 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3392 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3393 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3394 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3395 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3396 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3397 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3398 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3399 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3400 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3401 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3402 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3403 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3404 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3405 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3406 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3407 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3408 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3409 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3410 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3411 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3412 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3413 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3414 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3415 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3416 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3417 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3418 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3419 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3420 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3421 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3422 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3423 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3424 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3425 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3426 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3427 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3428 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3429 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3430 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3431 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3432 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3433 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3434 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3435 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3436 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3437 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3438 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3439 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3440 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3441 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3442 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3443 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3444 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3445 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3446 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3447 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3448 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3449 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3450 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3451 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3452 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3453 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3454 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3455 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3456 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3457 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3458 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3459 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3460 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3461 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3462 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3463 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3464 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3465 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3466 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3467 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3468 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3469 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3470 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3471 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3472 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3473 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3474 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3475 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3476 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3477 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3478 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3479 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3480 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3481 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3482 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3483 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3484 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3485 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3486 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3487 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3488 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3489 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3490 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3491 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3492 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3493 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3494 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3495 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3496 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3497 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3498 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3499 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3500 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3501 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3502 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3503 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3504 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3505 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3506 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3507 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3508 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3509 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3510 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3511 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3512 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3513 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3514 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3515 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3516 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3517 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3518 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3519 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3520 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3521 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3522 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3523 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3524 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3525 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3526 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3527 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3528 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3529 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3530 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3531 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3532 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3533 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3534 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3535 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3536 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3537 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3538 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3539 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3540 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3541 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3542 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3543 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3544 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3545 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3546 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3547 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3548 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3549 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3550 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3551 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3552 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3553 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3554 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3555 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3556 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3557 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3558 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3559 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3560 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3561 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3562 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3563 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3564 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3565 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3566 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3567 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3568 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3569 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3570 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3571 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3572 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3573 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3574 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3575 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3576 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3577 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3578 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3579 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3580 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3581 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3582 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3583 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3584 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3585 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3586 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3587 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3588 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3589 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3590 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3591 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3592 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3593 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3594 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3595 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3596 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3597 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3598 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3599 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3600 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3601 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3602 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3603 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3604 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3605 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3606 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3607 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3608 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3609 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3610 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3611 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3612 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3613 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3614 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3615 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3616 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3617 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3618 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3619 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3620 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3621 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3622 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3623 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3624 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3625 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3626 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3627 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3628 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3629 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3630 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3631 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3632 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3633 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3634 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3635 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3636 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3637 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3638 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3639 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3640 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3641 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3642 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3643 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3644 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3645 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3646 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3647 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3648 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3649 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3650 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3651 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3652 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3653 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3654 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3655 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3656 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3657 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3658 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3659 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3660 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3661 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3662 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3663 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3664 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3665 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3666 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3667 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3668 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3669 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3670 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3671 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3672 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3673 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3674 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3675 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3676 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3677 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3678 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3679 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3680 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3681 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3682 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3683 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3684 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3685 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3686 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3687 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3688 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3689 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3690 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3691 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3692 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3693 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3694 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3695 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3696 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3697 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3698 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3699 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3700 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3701 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3702 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3703 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3704 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3705 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3706 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3707 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3708 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3709 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3710 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3711 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3712 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3713 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3714 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3715 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3716 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3717 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3718 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3719 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3720 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3721 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3722 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3723 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3724 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3725 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3726 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3727 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3728 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3729 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3730 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3731 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3732 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3733 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3734 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3735 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3736 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3737 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3738 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3739 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3740 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3741 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3742 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3743 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3744 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3745 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3746 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3747 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3748 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3749 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3750 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3751 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3752 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3753 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3754 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3755 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3756 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3757 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3758 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3759 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3760 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3761 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3762 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3763 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3764 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3765 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3766 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3767 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3768 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3769 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3770 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3771 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3772 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3773 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3774 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3775 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3776 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3777 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3778 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3779 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3780 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3781 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3782 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3783 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3784 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3785 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3786 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3787 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3788 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3789 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3790 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3791 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3792 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3793 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3794 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3795 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3796 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3797 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3798 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3799 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3800 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3801 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3802 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3803 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3804 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3805 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3806 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3807 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3808 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3809 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3810 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3811 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3812 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3813 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3814 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3815 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3816 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3817 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3818 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3819 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3820 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3821 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3822 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3823 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3824 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3825 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3826 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3827 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3828 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3829 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3830 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3831 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3832 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3833 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3834 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3835 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3836 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3837 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3838 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3839 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3840 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3841 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3842 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3843 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3844 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3845 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3846 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3847 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3848 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3849 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3850 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3851 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3852 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3853 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3854 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3855 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3856 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3857 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3858 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3859 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3860 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3861 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3862 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3863 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3864 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3865 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3866 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3867 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3868 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3869 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3870 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3871 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3872 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3873 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3874 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3875 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3876 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3877 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3878 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3879 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3880 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3881 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3882 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3883 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3884 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3885 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3886 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3887 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3888 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3889 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3890 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3891 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3892 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3893 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3894 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3895 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3896 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3897 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3898 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3899 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3900 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3901 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3902 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3903 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3904 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3905 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3906 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3907 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3908 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3909 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3910 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3911 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3912 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3913 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3914 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3915 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3916 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3917 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3918 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3919 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3920 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3921 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3922 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3923 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3924 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3925 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3926 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3927 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3928 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3929 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3930 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3931 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3932 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3933 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3934 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3935 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3936 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3937 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3938 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3939 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3940 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3941 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3942 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3943 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3944 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3945 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3946 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3947 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3948 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3949 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3950 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3951 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3952 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3953 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3954 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3955 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3956 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3957 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3958 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3959 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3960 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3961 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3962 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3963 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3964 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3965 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3966 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3967 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3968 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3969 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3970 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3971 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3972 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3973 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3974 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3975 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3976 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3977 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3978 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3979 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3980 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3981 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3982 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3983 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3984 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3985 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3986 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3987 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3988 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3989 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3990 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3991 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3992 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3993 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3994 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3995 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3996 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3997 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3998 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3999 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4000 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4001 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4002 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4003 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4004 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4005 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4006 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4007 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4008 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4009 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4010 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4011 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4012 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4013 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4014 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4015 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4016 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4017 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4018 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4019 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4020 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4021 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4022 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4023 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4024 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4025 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4026 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4027 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4028 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4029 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4030 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4031 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4032 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4033 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4034 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4035 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4036 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4037 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4038 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4039 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4040 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4041 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4042 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4043 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4044 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4045 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4046 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4047 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4048 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4049 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4050 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4051 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4052 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4053 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4054 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4055 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4056 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4057 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4058 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4059 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4060 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4061 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4062 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4063 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4064 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4065 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4066 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4067 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4068 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4069 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4070 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4071 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4072 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4073 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4074 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4075 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4076 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4077 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4078 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4079 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4080 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4081 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4082 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4083 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4084 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4085 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4086 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4087 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4088 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4089 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4090 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4091 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4092 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4093 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4094 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4095 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4096 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4097 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4098 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4099 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4100 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4101 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4102 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4103 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4104 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4105 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4106 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4107 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4108 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4109 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4110 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4111 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4112 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4113 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4114 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4115 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4116 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4117 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4118 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4119 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4120 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4121 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4122 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4123 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4124 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4125 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4126 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4127 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4128 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4129 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4130 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4131 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4132 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4133 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4134 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4135 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4136 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4137 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4138 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4139 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4140 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4141 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4142 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4143 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4144 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4145 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4146 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4147 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4148 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4149 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4150 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4151 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4152 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4153 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4154 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4155 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4156 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4157 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4158 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4159 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4160 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4161 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4162 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4163 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4164 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4165 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4166 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4167 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4168 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4169 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4170 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4171 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4172 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4173 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4174 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4175 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4176 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4177 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4178 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4179 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4180 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4181 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4182 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4183 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4184 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4185 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4186 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4187 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4188 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4189 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4190 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4191 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4192 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4193 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4194 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4195 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4196 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4197 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4198 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4199 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4200 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4201 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4202 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4203 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4204 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4205 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4206 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4207 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4208 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4209 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4210 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4211 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4212 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4213 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4214 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4215 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4216 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4217 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4218 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4219 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4220 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4221 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4222 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4223 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4224 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4225 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4226 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4227 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4228 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4229 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4230 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4231 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4232 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4233 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4234 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4235 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4236 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4237 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4238 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4239 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4240 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4241 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4242 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4243 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4244 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4245 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4246 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4247 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4248 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4249 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4250 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4251 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4252 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4253 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4254 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4255 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4256 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4257 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4258 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4259 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4260 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4261 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4262 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4263 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4264 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4265 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4266 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4267 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4268 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4269 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4270 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4271 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4272 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4273 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4274 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4275 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4276 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4277 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4278 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4279 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4280 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4281 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4282 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4283 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4284 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4285 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4286 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4287 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4288 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4289 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4290 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4291 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4292 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4293 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4294 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4295 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4296 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4297 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4298 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4299 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4300 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4301 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4302 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4303 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4304 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4305 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4306 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4307 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4308 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4309 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4310 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4311 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4312 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4313 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4314 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4315 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4316 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4317 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4318 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4319 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4320 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4321 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4322 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4323 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4324 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4325 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4326 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4327 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4328 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4329 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4330 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4331 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4332 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4333 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4334 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4335 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4336 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4337 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4338 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4339 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4340 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4341 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4342 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4343 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4344 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4345 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4346 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4347 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4348 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4349 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4350 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4351 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4352 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4353 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4354 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4355 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4356 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4357 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4358 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4359 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4360 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4361 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4362 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4363 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4364 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4365 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4366 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4367 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4368 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4369 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4370 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4371 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4372 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4373 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4374 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4375 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4376 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4377 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4378 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4379 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4380 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4381 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4382 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4383 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4384 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4385 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4386 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4387 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4388 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4389 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4390 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4391 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4392 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4393 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4394 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4395 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4396 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4397 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4398 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4399 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4400 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4401 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4402 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4403 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4404 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4405 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4406 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4407 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4408 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4409 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4410 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4411 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4412 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4413 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4414 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4415 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4416 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4417 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4418 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4419 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4420 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4421 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4422 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4423 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4424 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4425 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4426 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4427 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4428 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4429 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4430 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4431 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4432 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4433 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4434 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4435 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4436 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4437 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4438 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4439 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4440 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4441 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4442 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4443 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4444 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4445 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4446 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4447 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4448 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4449 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4450 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4451 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4452 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4453 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4454 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4455 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4456 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4457 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4458 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4459 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4460 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4461 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4462 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4463 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4464 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4465 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4466 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4467 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4468 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4469 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4470 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4471 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4472 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4473 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4474 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4475 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4476 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4477 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4478 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4479 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4480 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4481 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4482 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4483 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4484 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4485 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4486 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4487 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4488 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4489 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4490 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4491 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4492 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4493 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4494 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4495 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4496 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4497 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4498 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4499 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4500 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4501 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4502 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4503 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4504 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4505 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4506 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4507 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4508 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4509 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4510 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4511 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4512 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4513 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4514 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4515 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4516 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4517 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4518 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4519 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4520 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4521 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4522 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4523 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4524 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4525 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4526 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4527 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4528 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4529 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4530 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4531 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4532 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4533 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4534 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4535 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4536 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4537 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4538 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4539 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4540 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4541 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4542 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4543 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4544 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4545 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4546 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4547 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4548 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4549 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4550 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4551 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4552 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4553 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4554 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4555 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4556 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4557 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4558 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4559 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4560 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4561 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4562 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4563 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4564 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4565 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4566 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4567 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4568 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4569 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4570 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4571 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4572 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4573 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4574 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4575 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4576 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4577 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4578 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4579 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4580 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4581 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4582 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4583 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4584 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4585 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4586 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4587 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4588 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4589 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4590 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4591 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4592 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4593 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4594 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4595 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4596 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4597 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4598 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4599 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4600 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4601 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4602 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4603 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4604 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4605 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4606 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4607 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4608 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4609 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4610 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4611 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4612 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4613 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4614 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4615 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4616 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4617 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4618 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4619 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4620 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4621 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4622 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4623 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4624 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4625 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4626 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4627 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4628 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4629 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4630 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4631 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4632 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4633 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4634 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4635 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4636 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4637 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4638 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4639 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4640 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4641 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4642 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4643 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4644 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4645 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4646 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4647 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4648 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4649 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4650 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4651 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4652 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4653 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4654 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4655 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4656 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4657 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4658 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4659 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4660 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4661 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4662 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4663 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4664 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4665 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4666 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4667 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4668 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4669 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4670 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4671 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4672 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4673 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4674 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4675 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4676 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4677 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4678 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4679 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4680 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4681 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4682 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4683 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4684 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4685 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4686 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4687 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4688 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4689 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4690 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4691 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4692 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4693 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4694 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4695 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4696 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4697 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4698 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4699 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4700 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4701 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4702 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4703 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4704 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4705 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4706 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4707 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4708 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4709 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4710 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4711 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4712 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4713 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4714 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4715 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4716 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4717 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4718 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4719 10bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4720 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4721 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4722 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4723 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4724 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4725 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4726 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4727 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4728 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4729 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4730 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4731 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4732 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4733 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4734 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4735 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4736 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4737 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4738 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4739 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d8 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4740 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4741 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4742 10bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4743 10bitdac_layout_0/9bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4744 10bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4745 10bitdac_layout_0/9bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4746 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4747 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4748 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d7 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4749 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4750 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4751 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4752 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4753 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4754 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4755 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4756 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4757 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4758 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4759 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4760 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4761 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4762 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4763 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4764 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4765 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4766 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4767 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4768 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4769 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4770 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4771 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4772 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4773 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4774 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4775 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4776 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4777 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4778 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4779 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4780 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4781 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4782 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4783 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4784 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4785 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4786 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4787 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4788 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4789 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4790 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4791 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4792 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4793 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4794 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4795 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4796 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4797 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4798 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4799 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4800 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4801 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4802 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4803 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4804 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4805 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4806 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4807 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4808 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4809 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4810 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4811 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4812 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4813 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4814 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4815 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4816 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4817 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4818 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4819 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4820 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4821 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4822 10bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4823 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4824 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4825 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4826 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4827 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4828 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4829 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4830 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4831 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4832 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4833 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4834 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4835 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4836 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4837 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4838 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4839 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4840 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4841 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4842 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4843 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4844 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4845 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4846 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4847 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4848 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4849 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4850 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4851 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4852 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4853 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4854 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4855 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4856 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4857 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4858 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4859 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4860 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4861 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4862 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4863 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4864 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4865 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4866 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4867 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4868 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4869 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4870 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4871 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4872 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4873 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4874 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4875 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4876 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4877 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4878 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4879 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4880 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4881 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4882 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4883 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4884 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4885 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4886 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4887 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4888 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4889 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4890 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4891 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4892 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4893 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4894 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4895 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4896 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4897 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4898 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4899 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4900 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4901 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4902 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4903 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4904 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4905 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4906 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4907 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4908 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4909 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4910 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4911 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4912 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4913 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4914 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4915 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4916 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4917 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4918 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4919 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4920 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4921 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4922 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4923 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4924 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4925 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4926 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4927 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4928 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4929 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4930 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4931 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4932 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4933 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4934 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4935 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4936 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4937 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4938 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4939 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4940 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4941 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4942 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4943 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4944 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4945 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4946 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4947 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4948 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4949 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4950 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4951 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4952 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4953 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4954 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4955 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4956 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4957 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4958 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4959 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4960 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4961 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4962 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4963 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4964 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4965 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4966 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4967 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4968 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4969 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4970 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4971 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4972 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4973 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4974 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4975 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4976 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4977 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4978 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4979 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4980 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4981 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4982 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4983 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4984 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4985 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4986 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4987 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4988 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4989 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4990 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4991 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4992 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4993 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4994 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4995 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4996 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4997 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4998 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4999 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5000 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5001 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5002 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5003 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5004 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5005 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5006 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5007 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5008 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5009 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5010 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5011 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5012 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5013 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5014 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5015 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5016 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5017 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5018 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5019 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5020 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5021 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5022 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5023 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5024 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5025 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5026 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5027 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5028 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5029 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5030 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5031 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5032 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5033 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5034 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5035 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5036 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5037 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5038 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5039 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5040 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5041 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5042 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5043 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5044 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5045 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5046 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5047 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5048 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5049 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5050 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5051 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5052 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5053 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5054 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5055 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5056 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5057 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5058 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5059 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5060 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5061 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5062 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5063 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5064 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5065 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5066 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5067 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5068 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5069 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5070 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5071 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5072 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5073 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5074 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5075 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5076 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5077 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5078 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5079 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5080 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5081 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5082 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5083 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5084 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5085 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5086 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5087 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5088 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5089 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5090 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5091 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5092 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5093 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5094 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5095 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5096 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5097 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5098 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5099 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5100 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5101 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5102 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5103 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5104 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5105 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5106 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5107 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5108 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5109 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5110 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5111 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5112 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5113 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5114 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5115 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5116 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5117 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5118 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5119 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5120 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5121 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5122 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5123 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5124 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5125 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5126 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5127 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5128 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5129 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5130 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5131 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5132 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5133 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5134 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5135 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5136 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5137 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5138 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5139 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5140 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5141 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5142 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5143 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5144 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5145 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5146 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5147 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5148 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5149 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5150 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5151 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5152 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5153 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5154 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5155 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5156 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5157 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5158 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5159 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5160 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5161 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5162 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5163 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5164 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5165 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5166 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5167 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5168 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5169 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5170 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5171 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5172 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5173 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5174 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5175 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5176 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5177 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5178 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5179 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5180 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5181 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5182 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5183 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5184 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5185 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5186 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5187 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5188 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5189 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5190 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5191 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5192 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5193 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5194 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5195 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5196 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5197 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5198 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5199 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5200 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5201 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5202 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5203 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5204 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5205 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5206 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5207 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5208 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5209 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5210 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5211 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5212 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5213 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5214 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5215 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5216 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5217 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5218 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5219 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5220 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5221 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5222 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5223 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5224 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5225 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5226 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5227 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5228 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5229 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5230 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5231 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5232 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5233 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5234 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5235 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5236 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5237 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5238 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5239 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5240 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5241 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5242 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5243 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5244 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5245 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5246 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5247 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5248 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5249 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5250 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5251 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5252 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5253 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5254 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5255 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5256 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5257 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5258 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5259 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5260 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5261 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5262 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5263 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5264 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5265 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5266 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5267 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5268 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5269 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5270 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5271 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5272 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5273 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5274 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5275 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5276 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5277 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5278 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5279 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5280 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5281 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5282 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5283 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5284 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5285 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5286 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5287 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5288 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5289 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5290 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5291 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5292 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5293 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5294 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5295 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5296 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5297 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5298 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5299 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5300 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5301 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5302 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5303 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5304 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5305 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5306 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5307 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5308 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5309 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5310 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5311 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5312 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5313 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5314 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5315 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5316 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5317 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5318 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5319 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5320 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5321 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5322 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5323 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5324 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5325 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5326 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5327 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5328 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5329 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5330 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5331 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5332 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5333 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5334 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5335 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5336 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5337 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5338 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5339 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5340 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5341 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5342 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5343 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5344 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5345 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5346 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5347 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5348 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5349 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5350 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5351 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5352 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5353 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5354 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5355 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5356 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5357 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5358 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5359 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5360 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5361 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5362 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5363 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5364 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5365 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5366 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5367 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5368 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5369 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5370 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5371 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5372 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5373 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5374 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5375 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5376 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5377 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5378 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5379 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5380 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5381 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5382 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5383 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5384 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5385 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5386 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5387 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5388 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5389 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5390 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5391 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5392 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5393 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5394 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5395 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5396 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5397 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5398 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5399 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5400 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5401 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5402 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5403 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5404 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5405 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5406 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5407 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5408 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5409 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5410 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5411 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5412 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5413 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5414 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5415 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5416 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5417 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5418 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5419 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5420 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5421 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5422 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5423 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5424 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5425 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5426 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5427 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5428 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5429 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5430 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5431 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5432 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5433 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5434 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5435 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5436 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5437 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5438 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5439 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5440 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5441 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5442 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5443 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5444 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5445 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5446 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5447 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5448 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5449 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5450 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5451 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5452 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5453 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5454 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5455 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5456 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5457 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5458 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5459 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5460 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5461 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5462 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5463 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5464 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5465 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5466 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5467 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5468 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5469 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5470 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5471 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5472 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5473 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5474 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5475 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5476 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5477 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5478 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5479 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5480 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5481 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5482 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5483 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5484 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5485 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5486 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5487 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5488 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5489 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5490 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5491 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5492 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5493 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5494 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5495 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5496 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5497 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5498 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5499 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5500 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5501 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5502 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5503 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5504 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5505 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5506 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5507 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5508 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5509 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5510 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5511 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5512 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5513 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5514 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5515 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5516 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5517 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5518 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5519 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5520 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5521 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5522 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5523 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5524 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5525 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5526 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5527 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5528 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5529 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5530 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5531 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5532 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5533 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5534 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5535 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5536 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5537 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5538 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5539 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5540 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5541 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5542 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5543 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5544 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5545 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5546 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5547 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5548 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5549 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5550 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5551 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5552 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5553 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5554 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5555 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5556 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5557 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5558 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5559 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5560 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5561 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5562 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5563 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5564 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5565 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5566 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5567 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5568 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5569 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5570 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5571 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5572 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5573 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5574 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5575 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5576 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5577 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5578 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5579 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5580 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5581 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5582 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5583 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5584 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5585 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5586 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5587 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5588 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5589 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5590 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5591 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5592 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5593 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5594 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5595 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5596 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5597 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5598 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5599 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5600 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5601 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5602 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5603 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5604 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5605 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5606 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5607 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5608 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5609 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5610 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5611 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5612 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5613 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5614 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5615 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5616 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5617 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5618 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5619 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5620 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5621 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5622 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5623 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5624 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5625 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5626 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5627 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5628 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5629 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5630 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5631 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5632 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5633 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5634 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5635 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5636 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5637 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5638 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5639 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5640 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5641 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5642 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5643 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5644 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5645 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5646 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5647 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5648 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5649 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5650 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5651 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5652 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5653 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5654 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5655 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5656 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5657 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5658 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5659 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5660 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5661 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5662 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5663 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5664 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5665 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5666 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5667 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5668 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5669 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5670 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5671 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5672 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5673 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5674 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5675 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5676 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5677 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5678 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5679 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5680 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5681 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5682 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5683 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5684 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5685 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5686 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5687 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5688 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5689 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5690 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5691 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5692 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5693 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5694 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5695 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5696 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5697 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5698 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5699 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5700 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5701 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5702 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5703 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5704 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5705 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5706 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5707 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5708 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5709 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5710 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5711 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5712 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5713 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5714 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5715 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5716 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5717 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5718 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5719 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5720 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5721 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5722 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5723 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5724 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5725 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5726 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5727 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5728 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5729 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5730 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5731 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5732 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5733 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5734 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5735 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5736 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5737 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5738 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5739 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5740 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5741 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5742 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5743 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5744 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5745 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5746 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5747 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5748 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5749 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5750 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5751 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5752 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5753 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5754 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5755 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5756 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5757 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5758 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5759 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5760 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5761 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5762 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5763 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5764 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5765 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5766 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5767 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5768 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5769 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5770 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5771 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5772 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5773 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5774 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5775 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5776 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5777 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5778 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5779 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5780 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5781 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5782 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5783 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5784 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5785 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5786 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5787 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5788 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5789 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5790 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5791 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5792 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5793 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5794 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5795 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5796 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5797 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5798 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5799 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5800 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5801 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5802 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5803 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5804 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5805 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5806 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5807 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5808 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5809 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5810 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5811 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5812 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5813 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5814 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5815 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5816 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5817 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5818 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5819 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5820 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5821 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5822 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5823 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5824 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5825 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5826 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5827 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5828 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5829 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5830 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5831 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5832 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5833 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5834 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5835 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5836 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5837 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5838 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5839 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5840 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5841 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5842 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5843 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5844 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5845 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5846 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5847 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5848 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5849 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5850 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5851 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5852 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5853 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5854 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5855 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5856 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5857 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5858 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5859 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5860 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5861 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5862 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5863 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5864 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5865 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5866 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5867 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5868 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5869 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5870 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5871 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5872 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5873 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5874 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5875 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5876 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5877 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5878 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5879 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5880 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5881 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5882 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5883 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5884 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5885 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5886 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5887 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5888 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5889 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5890 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5891 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5892 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5893 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5894 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5895 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5896 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5897 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5898 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5899 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5900 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5901 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5902 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5903 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5904 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5905 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5906 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5907 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5908 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5909 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5910 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5911 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5912 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5913 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5914 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5915 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5916 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5917 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5918 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5919 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5920 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5921 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5922 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5923 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5924 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5925 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5926 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5927 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5928 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5929 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5930 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5931 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5932 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5933 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5934 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5935 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5936 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5937 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5938 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5939 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5940 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5941 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5942 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5943 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5944 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5945 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5946 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5947 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5948 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5949 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5950 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5951 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5952 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5953 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5954 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5955 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5956 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5957 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5958 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5959 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5960 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5961 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5962 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5963 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5964 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5965 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5966 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5967 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5968 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5969 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5970 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5971 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5972 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5973 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5974 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5975 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5976 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5977 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5978 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5979 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5980 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5981 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5982 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5983 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5984 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5985 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5986 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5987 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5988 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5989 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5990 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5991 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5992 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5993 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5994 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5995 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5996 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5997 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5998 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5999 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6000 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6001 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6002 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6003 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6004 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6005 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6006 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6007 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6008 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6009 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6010 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6011 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6012 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6013 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6014 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6015 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6016 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6017 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6018 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6019 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6020 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6021 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6022 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6023 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6024 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6025 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6026 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6027 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6028 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6029 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6030 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6031 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6032 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6033 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6034 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6035 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6036 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6037 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6038 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6039 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6040 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6041 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6042 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6043 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6044 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6045 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6046 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6047 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6048 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6049 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6050 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6051 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6052 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6053 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6054 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6055 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6056 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6057 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6058 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6059 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6060 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6061 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6062 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6063 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6064 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6065 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6066 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6067 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6068 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6069 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6070 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6071 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6072 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6073 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6074 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6075 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6076 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6077 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6078 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6079 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6080 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6081 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6082 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6083 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6084 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6085 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6086 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6087 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6088 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6089 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6090 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6091 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6092 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6093 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6094 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6095 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6096 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6097 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6098 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6099 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6100 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6101 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6102 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6103 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6104 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6105 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6106 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6107 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6108 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6109 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6110 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6111 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6112 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6113 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6114 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6115 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6116 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6117 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6118 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6119 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6120 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6121 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6122 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6123 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6124 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6125 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6126 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6127 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6128 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6129 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6130 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6131 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6132 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6133 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6134 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6135 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6136 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6137 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6138 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6139 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6140 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6141 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6142 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6143 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6144 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6145 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6146 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6147 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6148 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6149 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6150 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6151 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6152 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6153 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6154 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6155 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6156 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6157 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6158 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6159 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6160 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6161 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6162 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6163 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6164 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6165 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6166 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6167 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6168 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6169 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6170 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6171 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6172 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6173 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6174 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6175 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6176 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6177 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6178 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6179 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6180 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6181 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6182 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6183 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6184 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6185 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6186 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6187 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6188 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6189 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6190 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6191 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6192 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6193 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6194 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6195 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6196 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6197 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6198 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6199 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6200 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6201 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6202 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6203 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6204 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6205 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6206 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6207 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6208 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6209 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6210 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6211 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6212 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6213 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6214 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6215 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6216 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6217 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6218 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6219 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6220 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6221 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6222 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6223 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6224 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6225 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6226 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6227 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6228 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6229 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6230 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6231 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6232 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6233 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6234 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6235 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6236 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6237 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6238 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6239 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6240 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6241 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6242 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6243 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6244 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6245 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6246 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6247 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6248 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6249 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6250 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6251 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6252 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6253 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6254 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6255 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6256 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6257 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6258 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6259 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6260 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6261 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6262 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6263 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6264 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6265 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6266 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6267 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6268 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6269 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6270 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6271 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6272 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6273 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6274 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6275 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6276 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6277 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6278 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6279 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6280 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6281 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6282 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6283 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6284 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6285 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6286 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6287 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6288 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6289 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6290 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6291 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6292 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6293 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6294 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6295 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6296 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6297 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6298 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6299 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6300 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6301 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6302 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6303 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6304 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6305 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6306 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6307 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6308 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6309 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6310 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6311 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6312 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6313 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6314 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6315 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6316 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6317 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6318 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6319 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6320 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6321 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6322 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6323 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6324 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6325 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6326 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6327 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6328 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6329 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6330 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6331 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6332 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6333 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6334 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6335 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6336 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6337 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6338 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6339 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6340 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6341 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6342 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6343 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6344 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6345 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6346 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6347 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6348 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6349 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6350 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6351 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6352 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6353 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6354 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6355 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6356 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6357 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6358 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6359 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6360 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6361 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6362 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6363 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6364 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6365 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6366 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6367 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6368 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6369 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6370 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6371 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6372 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6373 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6374 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6375 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6376 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6377 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6378 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6379 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6380 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6381 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6382 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6383 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6384 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6385 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6386 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6387 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6388 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6389 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6390 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6391 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6392 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6393 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6394 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6395 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6396 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6397 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6398 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6399 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6400 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6401 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6402 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6403 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6404 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6405 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6406 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6407 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6408 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6409 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6410 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6411 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6412 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6413 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6414 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6415 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6416 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6417 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6418 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6419 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6420 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6421 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6422 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6423 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6424 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6425 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6426 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6427 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6428 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6429 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6430 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6431 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6432 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6433 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6434 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6435 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6436 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6437 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6438 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6439 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6440 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6441 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6442 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6443 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6444 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6445 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6446 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6447 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6448 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6449 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6450 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6451 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6452 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6453 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6454 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6455 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6456 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6457 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6458 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6459 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6460 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6461 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6462 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6463 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6464 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6465 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6466 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6467 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6468 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6469 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6470 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6471 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6472 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6473 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6474 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6475 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6476 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6477 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6478 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6479 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6480 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6481 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6482 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6483 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6484 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6485 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6486 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6487 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6488 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6489 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6490 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6491 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6492 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6493 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6494 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6495 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6496 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6497 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6498 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6499 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6500 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6501 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6502 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6503 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6504 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6505 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6506 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6507 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6508 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6509 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6510 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6511 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6512 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6513 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6514 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6515 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6516 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6517 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6518 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6519 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6520 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6521 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6522 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6523 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6524 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6525 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6526 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6527 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6528 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6529 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6530 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6531 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6532 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6533 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6534 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6535 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6536 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6537 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6538 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6539 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6540 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6541 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6542 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6543 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6544 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6545 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6546 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6547 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6548 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6549 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6550 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6551 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6552 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6553 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6554 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6555 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6556 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6557 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6558 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6559 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6560 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6561 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6562 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6563 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6564 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6565 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6566 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6567 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6568 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6569 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6570 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6571 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6572 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6573 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6574 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6575 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6576 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6577 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6578 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6579 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6580 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6581 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6582 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6583 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6584 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6585 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6586 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6587 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6588 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6589 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6590 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6591 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6592 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6593 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6594 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6595 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6596 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6597 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6598 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6599 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6600 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6601 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6602 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6603 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6604 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6605 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6606 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6607 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6608 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6609 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6610 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6611 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6612 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6613 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6614 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6615 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6616 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6617 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6618 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6619 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6620 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6621 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6622 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6623 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6624 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6625 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6626 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6627 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6628 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6629 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6630 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6631 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6632 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6633 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6634 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6635 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6636 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6637 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6638 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6639 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6640 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6641 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6642 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6643 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6644 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6645 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6646 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6647 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6648 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6649 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6650 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6651 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6652 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6653 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6654 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6655 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6656 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6657 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6658 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6659 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6660 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6661 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6662 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6663 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6664 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6665 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6666 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6667 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6668 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6669 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6670 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6671 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6672 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6673 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6674 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6675 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6676 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6677 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6678 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6679 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6680 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6681 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6682 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6683 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6684 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6685 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6686 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6687 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6688 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6689 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6690 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6691 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6692 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6693 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6694 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6695 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6696 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6697 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6698 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6699 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6700 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6701 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6702 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6703 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6704 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6705 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6706 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6707 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6708 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6709 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6710 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6711 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6712 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6713 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6714 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6715 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6716 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6717 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6718 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6719 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6720 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6721 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6722 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6723 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6724 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6725 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6726 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6727 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6728 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6729 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6730 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6731 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6732 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6733 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6734 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6735 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6736 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6737 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6738 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6739 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6740 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6741 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6742 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6743 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6744 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6745 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6746 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6747 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6748 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6749 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6750 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6751 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6752 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6753 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6754 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6755 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6756 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6757 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6758 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6759 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6760 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6761 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6762 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6763 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6764 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6765 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6766 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6767 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6768 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6769 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6770 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6771 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6772 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6773 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6774 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6775 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6776 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6777 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6778 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6779 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6780 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6781 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6782 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6783 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6784 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6785 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6786 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6787 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6788 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6789 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6790 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6791 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6792 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6793 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6794 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6795 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6796 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6797 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6798 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6799 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6800 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6801 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6802 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6803 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6804 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6805 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6806 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6807 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6808 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6809 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6810 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6811 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6812 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6813 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6814 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6815 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6816 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6817 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6818 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6819 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6820 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6821 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6822 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6823 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6824 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6825 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6826 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6827 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6828 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6829 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6830 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6831 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6832 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6833 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6834 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6835 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6836 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6837 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6838 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6839 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6840 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6841 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6842 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6843 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6844 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6845 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6846 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6847 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6848 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6849 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6850 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6851 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6852 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6853 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6854 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6855 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6856 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6857 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6858 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6859 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6860 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6861 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6862 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6863 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6864 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6865 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6866 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6867 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6868 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6869 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6870 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6871 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6872 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6873 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6874 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6875 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6876 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6877 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6878 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6879 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6880 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6881 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6882 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6883 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6884 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6885 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6886 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6887 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6888 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6889 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6890 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6891 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6892 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6893 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6894 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6895 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6896 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6897 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6898 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6899 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6900 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6901 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6902 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6903 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6904 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6905 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6906 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6907 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6908 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6909 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6910 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6911 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6912 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6913 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6914 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6915 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6916 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6917 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6918 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6919 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6920 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6921 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6922 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6923 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6924 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6925 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6926 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6927 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6928 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6929 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6930 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6931 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6932 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6933 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6934 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6935 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6936 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6937 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6938 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6939 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6940 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6941 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6942 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6943 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6944 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6945 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6946 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6947 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6948 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6949 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6950 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6951 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6952 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6953 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6954 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6955 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6956 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6957 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6958 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6959 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6960 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6961 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6962 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6963 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6964 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6965 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6966 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6967 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6968 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6969 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6970 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6971 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6972 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6973 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6974 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6975 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6976 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6977 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6978 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6979 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6980 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6981 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6982 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6983 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6984 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6985 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6986 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6987 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6988 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6989 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6990 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6991 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6992 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6993 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6994 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6995 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6996 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6997 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6998 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6999 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7000 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7001 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7002 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7003 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7004 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7005 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7006 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7007 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7008 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7009 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7010 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7011 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7012 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7013 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7014 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7015 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7016 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7017 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7018 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7019 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7020 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7021 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7022 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7023 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7024 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7025 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7026 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7027 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7028 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7029 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7030 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7031 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7032 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7033 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7034 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7035 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7036 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7037 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7038 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7039 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7040 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7041 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7042 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7043 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7044 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7045 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7046 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7047 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7048 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7049 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7050 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7051 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7052 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7053 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7054 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7055 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7056 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7057 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7058 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7059 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7060 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7061 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7062 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7063 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7064 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7065 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7066 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7067 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7068 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7069 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7070 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7071 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7072 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7073 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7074 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7075 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7076 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7077 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7078 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7079 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7080 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7081 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7082 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7083 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7084 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7085 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7086 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7087 10bitdac_layout_0/9bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7088 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7089 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7090 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7091 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7092 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7093 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7094 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7095 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7096 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7097 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7098 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7099 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7100 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7101 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7102 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7103 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7104 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7105 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7106 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7107 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d7 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7108 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7109 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7110 10bitdac_layout_0/9bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7111 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7112 10bitdac_layout_0/9bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7113 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7114 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7115 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7116 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7117 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7118 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7119 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7120 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7121 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7122 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7123 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7124 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7125 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7126 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7127 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7128 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7129 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7130 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7131 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7132 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7133 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7134 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7135 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7136 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7137 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7138 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7139 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7140 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7141 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7142 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7143 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7144 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7145 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7146 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7147 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7148 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7149 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7150 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7151 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7152 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7153 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7154 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7155 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7156 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7157 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7158 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7159 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7160 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7161 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7162 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7163 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7164 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7165 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7166 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7167 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7168 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7169 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7170 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7171 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7172 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7173 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7174 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7175 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7176 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7177 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7178 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7179 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7180 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7181 10bitdac_layout_0/9bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7182 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7183 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7184 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7185 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7186 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7187 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7188 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7189 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7190 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7191 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7192 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7193 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7194 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7195 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7196 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7197 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7198 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7199 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7200 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7201 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7202 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7203 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7204 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7205 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7206 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7207 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7208 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7209 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7210 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7211 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7212 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7213 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7214 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7215 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7216 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7217 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7218 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7219 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7220 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7221 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7222 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7223 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7224 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7225 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7226 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7227 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7228 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7229 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7230 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7231 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7232 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7233 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7234 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7235 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7236 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7237 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7238 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7239 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7240 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7241 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7242 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7243 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7244 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7245 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7246 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7247 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7248 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7249 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7250 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7251 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7252 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7253 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7254 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7255 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7256 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7257 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7258 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7259 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7260 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7261 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7262 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7263 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7264 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7265 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7266 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7267 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7268 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7269 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7270 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7271 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7272 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7273 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7274 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7275 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7276 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7277 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7278 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7279 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7280 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7281 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7282 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7283 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7284 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7285 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7286 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7287 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7288 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7289 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7290 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7291 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7292 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7293 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7294 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7295 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7296 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7297 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7298 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7299 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7300 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7301 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7302 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7303 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7304 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7305 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7306 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7307 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7308 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7309 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7310 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7311 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7312 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7313 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7314 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7315 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7316 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7317 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7318 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7319 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7320 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7321 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7322 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7323 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7324 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7325 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7326 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7327 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7328 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7329 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7330 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7331 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7332 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7333 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7334 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7335 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7336 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7337 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7338 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7339 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7340 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7341 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7342 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7343 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7344 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7345 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7346 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7347 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7348 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7349 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7350 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7351 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7352 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7353 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7354 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7355 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7356 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7357 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7358 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7359 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7360 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7361 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7362 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7363 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7364 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7365 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7366 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7367 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7368 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7369 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7370 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7371 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7372 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7373 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7374 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7375 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7376 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7377 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7378 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7379 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7380 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7381 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7382 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7383 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7384 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7385 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7386 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7387 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7388 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7389 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7390 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7391 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7392 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7393 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7394 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7395 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7396 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7397 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7398 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7399 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7400 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7401 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7402 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7403 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7404 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7405 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7406 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7407 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7408 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7409 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7410 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7411 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7412 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7413 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7414 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7415 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7416 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7417 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7418 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7419 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7420 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7421 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7422 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7423 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7424 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7425 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7426 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7427 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7428 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7429 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7430 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7431 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7432 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7433 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7434 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7435 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7436 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7437 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7438 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7439 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7440 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7441 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7442 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7443 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7444 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7445 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7446 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7447 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7448 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7449 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7450 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7451 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7452 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7453 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7454 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7455 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7456 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7457 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7458 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7459 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7460 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7461 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7462 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7463 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7464 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7465 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7466 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7467 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7468 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7469 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7470 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7471 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7472 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7473 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7474 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7475 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7476 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7477 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7478 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7479 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7480 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7481 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7482 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7483 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7484 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7485 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7486 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7487 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7488 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7489 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7490 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7491 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7492 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7493 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7494 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7495 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7496 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7497 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7498 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7499 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7500 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7501 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7502 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7503 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7504 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7505 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7506 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7507 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7508 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7509 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7510 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7511 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7512 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7513 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7514 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7515 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7516 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7517 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7518 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7519 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7520 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7521 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7522 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7523 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7524 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7525 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7526 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7527 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7528 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7529 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7530 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7531 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7532 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7533 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7534 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7535 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7536 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7537 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7538 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7539 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7540 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7541 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7542 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7543 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7544 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7545 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7546 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7547 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7548 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7549 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7550 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7551 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7552 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7553 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7554 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7555 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7556 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7557 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7558 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7559 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7560 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7561 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7562 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7563 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7564 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7565 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7566 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7567 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7568 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7569 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7570 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7571 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7572 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7573 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7574 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7575 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7576 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7577 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7578 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7579 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7580 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7581 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7582 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7583 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7584 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7585 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7586 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7587 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7588 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7589 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7590 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7591 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7592 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7593 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7594 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7595 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7596 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7597 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7598 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7599 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7600 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7601 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7602 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7603 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7604 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7605 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7606 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7607 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7608 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7609 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7610 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7611 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7612 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7613 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7614 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7615 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7616 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7617 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7618 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7619 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7620 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7621 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7622 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7623 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7624 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7625 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7626 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7627 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7628 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7629 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7630 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7631 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7632 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7633 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7634 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7635 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7636 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7637 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7638 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7639 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7640 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7641 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7642 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7643 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7644 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7645 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7646 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7647 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7648 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7649 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7650 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7651 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7652 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7653 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7654 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7655 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7656 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7657 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7658 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7659 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7660 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7661 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7662 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7663 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7664 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7665 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7666 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7667 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7668 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7669 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7670 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7671 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7672 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7673 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7674 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7675 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7676 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7677 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7678 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7679 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7680 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7681 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7682 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7683 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7684 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7685 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7686 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7687 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7688 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7689 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7690 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7691 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7692 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7693 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7694 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7695 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7696 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7697 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7698 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7699 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7700 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7701 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7702 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7703 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7704 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7705 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7706 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7707 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7708 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7709 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7710 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7711 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7712 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7713 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7714 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7715 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7716 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7717 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7718 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7719 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7720 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7721 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7722 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7723 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7724 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7725 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7726 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7727 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7728 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7729 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7730 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7731 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7732 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7733 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7734 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7735 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7736 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7737 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7738 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7739 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7740 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7741 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7742 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7743 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7744 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7745 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7746 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7747 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7748 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7749 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7750 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7751 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7752 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7753 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7754 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7755 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7756 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7757 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7758 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7759 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7760 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7761 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7762 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7763 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7764 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7765 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7766 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7767 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7768 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7769 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7770 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7771 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7772 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7773 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7774 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7775 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7776 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7777 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7778 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7779 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7780 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7781 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7782 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7783 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7784 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7785 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7786 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7787 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7788 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7789 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7790 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7791 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7792 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7793 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7794 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7795 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7796 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7797 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7798 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7799 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7800 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7801 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7802 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7803 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7804 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7805 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7806 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7807 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7808 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7809 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7810 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7811 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7812 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7813 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7814 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7815 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7816 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7817 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7818 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7819 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7820 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7821 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7822 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7823 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7824 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7825 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7826 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7827 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7828 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7829 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7830 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7831 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7832 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7833 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7834 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7835 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7836 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7837 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7838 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7839 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7840 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7841 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7842 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7843 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7844 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7845 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7846 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7847 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7848 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7849 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7850 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7851 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7852 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7853 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7854 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7855 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7856 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7857 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7858 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7859 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7860 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7861 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7862 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7863 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7864 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7865 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7866 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7867 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7868 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7869 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7870 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7871 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7872 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7873 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7874 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7875 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7876 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7877 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7878 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7879 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7880 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7881 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7882 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7883 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7884 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7885 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7886 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7887 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7888 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7889 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7890 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7891 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7892 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7893 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7894 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7895 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7896 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7897 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7898 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7899 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7900 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7901 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7902 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7903 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7904 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7905 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7906 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7907 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7908 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7909 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7910 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7911 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7912 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7913 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7914 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7915 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7916 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7917 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7918 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7919 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7920 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7921 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7922 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7923 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7924 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7925 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7926 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7927 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7928 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7929 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7930 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7931 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7932 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7933 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7934 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7935 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7936 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7937 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7938 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7939 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7940 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7941 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7942 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7943 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7944 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7945 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7946 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7947 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7948 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7949 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7950 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7951 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7952 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7953 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7954 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7955 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7956 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7957 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7958 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7959 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7960 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7961 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7962 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7963 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7964 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7965 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7966 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7967 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7968 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7969 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7970 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7971 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7972 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7973 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7974 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7975 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7976 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7977 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7978 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7979 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7980 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7981 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7982 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7983 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7984 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7985 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7986 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7987 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7988 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7989 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7990 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7991 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7992 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7993 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7994 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7995 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7996 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7997 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7998 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7999 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8000 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8001 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8002 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8003 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8004 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8005 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8006 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8007 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8008 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8009 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8010 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8011 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8012 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8013 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8014 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8015 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8016 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8017 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8018 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8019 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8020 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8021 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8022 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8023 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8024 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8025 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8026 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8027 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8028 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8029 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8030 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8031 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8032 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8033 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8034 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8035 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8036 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8037 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8038 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8039 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8040 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8041 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8042 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8043 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8044 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8045 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8046 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8047 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8048 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8049 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8050 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8051 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8052 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8053 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8054 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8055 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8056 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8057 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8058 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8059 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8060 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8061 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8062 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8063 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8064 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8065 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8066 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8067 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8068 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8069 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8070 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8071 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8072 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8073 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8074 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8075 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8076 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8077 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8078 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8079 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8080 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8081 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8082 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8083 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8084 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8085 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8086 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8087 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8088 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8089 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8090 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8091 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8092 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8093 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8094 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8095 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8096 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8097 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8098 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8099 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8100 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8101 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8102 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8103 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8104 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8105 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8106 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8107 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8108 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8109 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8110 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8111 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8112 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8113 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8114 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8115 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8116 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8117 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8118 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8119 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8120 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8121 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8122 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8123 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8124 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8125 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8126 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8127 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8128 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8129 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8130 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8131 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8132 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8133 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8134 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8135 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8136 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8137 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8138 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8139 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8140 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8141 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8142 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8143 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8144 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8145 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8146 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8147 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8148 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8149 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8150 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8151 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8152 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8153 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8154 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8155 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8156 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8157 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8158 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8159 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8160 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8161 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8162 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8163 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8164 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8165 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8166 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8167 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8168 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8169 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8170 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8171 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8172 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8173 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8174 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8175 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8176 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8177 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8178 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8179 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8180 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8181 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8182 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8183 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8184 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8185 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8186 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8187 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8188 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8189 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8190 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8191 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8192 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8193 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8194 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8195 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8196 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8197 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8198 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8199 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8200 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8201 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8202 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8203 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8204 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8205 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8206 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8207 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8208 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8209 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8210 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8211 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8212 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8213 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8214 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8215 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8216 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8217 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8218 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8219 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8220 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8221 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8222 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8223 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8224 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8225 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8226 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8227 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8228 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8229 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8230 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8231 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8232 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8233 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8234 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8235 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8236 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8237 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8238 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8239 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8240 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8241 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8242 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8243 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8244 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8245 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8246 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8247 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8248 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8249 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8250 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8251 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8252 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8253 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8254 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8255 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8256 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8257 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8258 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8259 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8260 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8261 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8262 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8263 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8264 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8265 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8266 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8267 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8268 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8269 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8270 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8271 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8272 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8273 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8274 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8275 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8276 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8277 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8278 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8279 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8280 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8281 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8282 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8283 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8284 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8285 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8286 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8287 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8288 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8289 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8290 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8291 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8292 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8293 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8294 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8295 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8296 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8297 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8298 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8299 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8300 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8301 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8302 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8303 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8304 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8305 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8306 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8307 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8308 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8309 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8310 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8311 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8312 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8313 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8314 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8315 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8316 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8317 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8318 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8319 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8320 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8321 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8322 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8323 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8324 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8325 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8326 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8327 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8328 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8329 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8330 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8331 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8332 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8333 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8334 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8335 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8336 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8337 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8338 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8339 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8340 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8341 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8342 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8343 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8344 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8345 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8346 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8347 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8348 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8349 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8350 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8351 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8352 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8353 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8354 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8355 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8356 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8357 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8358 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8359 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8360 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8361 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8362 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8363 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8364 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8365 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8366 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8367 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8368 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8369 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8370 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8371 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8372 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8373 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8374 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8375 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8376 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8377 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8378 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8379 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8380 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8381 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8382 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8383 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8384 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8385 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8386 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8387 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8388 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8389 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8390 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8391 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8392 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8393 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8394 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8395 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8396 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8397 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8398 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8399 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8400 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8401 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8402 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8403 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8404 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8405 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8406 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8407 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8408 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8409 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8410 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8411 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8412 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8413 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8414 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8415 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8416 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8417 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8418 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8419 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8420 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8421 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8422 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8423 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8424 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8425 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8426 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8427 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8428 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8429 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8430 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8431 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8432 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8433 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8434 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8435 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8436 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8437 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8438 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8439 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8440 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8441 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8442 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8443 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8444 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8445 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8446 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8447 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8448 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8449 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8450 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8451 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8452 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8453 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8454 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8455 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8456 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8457 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8458 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8459 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8460 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8461 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8462 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8463 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8464 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8465 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8466 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8467 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8468 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8469 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8470 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8471 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8472 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8473 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8474 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8475 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8476 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8477 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8478 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8479 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8480 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8481 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8482 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8483 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8484 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8485 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8486 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8487 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8488 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8489 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8490 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8491 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8492 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8493 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8494 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8495 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8496 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8497 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8498 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8499 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8500 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8501 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8502 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8503 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8504 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8505 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8506 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8507 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8508 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8509 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8510 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8511 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8512 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8513 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8514 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8515 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8516 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8517 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8518 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8519 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8520 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8521 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8522 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8523 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8524 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8525 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8526 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8527 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8528 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8529 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8530 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8531 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8532 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8533 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8534 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8535 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8536 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8537 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8538 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8539 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8540 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8541 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8542 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8543 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8544 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8545 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8546 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8547 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8548 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8549 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8550 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8551 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8552 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8553 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8554 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8555 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8556 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8557 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8558 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8559 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8560 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8561 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8562 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8563 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8564 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8565 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8566 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8567 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8568 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8569 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8570 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8571 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8572 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8573 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8574 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8575 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8576 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8577 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8578 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8579 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8580 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8581 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8582 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8583 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8584 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8585 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8586 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8587 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8588 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8589 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8590 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8591 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8592 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8593 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8594 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8595 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8596 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8597 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8598 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8599 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8600 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8601 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8602 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8603 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8604 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8605 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8606 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8607 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8608 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8609 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8610 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8611 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8612 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8613 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8614 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8615 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8616 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8617 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8618 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8619 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8620 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8621 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8622 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8623 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8624 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8625 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8626 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8627 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8628 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8629 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8630 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8631 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8632 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8633 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8634 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8635 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8636 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8637 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8638 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8639 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8640 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8641 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8642 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8643 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8644 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8645 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8646 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8647 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8648 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8649 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8650 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8651 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8652 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8653 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8654 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8655 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8656 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8657 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8658 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8659 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8660 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8661 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8662 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8663 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8664 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8665 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8666 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8667 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8668 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8669 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8670 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8671 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8672 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8673 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8674 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8675 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8676 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8677 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8678 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8679 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8680 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8681 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8682 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8683 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8684 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8685 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8686 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8687 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8688 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8689 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8690 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8691 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8692 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8693 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8694 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8695 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8696 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8697 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8698 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8699 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8700 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8701 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8702 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8703 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8704 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8705 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8706 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8707 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8708 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8709 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8710 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8711 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8712 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8713 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8714 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8715 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8716 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8717 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8718 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8719 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8720 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8721 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8722 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8723 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8724 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8725 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8726 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8727 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8728 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8729 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8730 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8731 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8732 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8733 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8734 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8735 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8736 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8737 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8738 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8739 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8740 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8741 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8742 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8743 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8744 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8745 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8746 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8747 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8748 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8749 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8750 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8751 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8752 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8753 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8754 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8755 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8756 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8757 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8758 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8759 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8760 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8761 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8762 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8763 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8764 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8765 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8766 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8767 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8768 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8769 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8770 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8771 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8772 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8773 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8774 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8775 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8776 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8777 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8778 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8779 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8780 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8781 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8782 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8783 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8784 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8785 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8786 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8787 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8788 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8789 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8790 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8791 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8792 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8793 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8794 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8795 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8796 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8797 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8798 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8799 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8800 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8801 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8802 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8803 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8804 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8805 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8806 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8807 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8808 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8809 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8810 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8811 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8812 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8813 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8814 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8815 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8816 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8817 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8818 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8819 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8820 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8821 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8822 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8823 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8824 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8825 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8826 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8827 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8828 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8829 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8830 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8831 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8832 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8833 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8834 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8835 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8836 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8837 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8838 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8839 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8840 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8841 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8842 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8843 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8844 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8845 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8846 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8847 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8848 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8849 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8850 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8851 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8852 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8853 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8854 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8855 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8856 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8857 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8858 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8859 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8860 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8861 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8862 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8863 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8864 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8865 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8866 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8867 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8868 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8869 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8870 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8871 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8872 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8873 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8874 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8875 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8876 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8877 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8878 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8879 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8880 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8881 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8882 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8883 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8884 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8885 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8886 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8887 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8888 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8889 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8890 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8891 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8892 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8893 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8894 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8895 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8896 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8897 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8898 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8899 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8900 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8901 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8902 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8903 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8904 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8905 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8906 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8907 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8908 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8909 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8910 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8911 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8912 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8913 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8914 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8915 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8916 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8917 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8918 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8919 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8920 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8921 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8922 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8923 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8924 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8925 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8926 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8927 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8928 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8929 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8930 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8931 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8932 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8933 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8934 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8935 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8936 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8937 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8938 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8939 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8940 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8941 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8942 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8943 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8944 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8945 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8946 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8947 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8948 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8949 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8950 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8951 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8952 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8953 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8954 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8955 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8956 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8957 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8958 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8959 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8960 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8961 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8962 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8963 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8964 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8965 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8966 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8967 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8968 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8969 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8970 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8971 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8972 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8973 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8974 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8975 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8976 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8977 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8978 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8979 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8980 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8981 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8982 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8983 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8984 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8985 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8986 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8987 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8988 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8989 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8990 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8991 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8992 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8993 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8994 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8995 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8996 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8997 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8998 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8999 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9000 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9001 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9002 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9003 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9004 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9005 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9006 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9007 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9008 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9009 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9010 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9011 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9012 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9013 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9014 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9015 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9016 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9017 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9018 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9019 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9020 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9021 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9022 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9023 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9024 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9025 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9026 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9027 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9028 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9029 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9030 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9031 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9032 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9033 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9034 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9035 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9036 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9037 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9038 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9039 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9040 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9041 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9042 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9043 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9044 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9045 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9046 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9047 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9048 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9049 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9050 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9051 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9052 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9053 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9054 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9055 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9056 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9057 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9058 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9059 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9060 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9061 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9062 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9063 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9064 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9065 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9066 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9067 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9068 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9069 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9070 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9071 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9072 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9073 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9074 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9075 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9076 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9077 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9078 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9079 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9080 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9081 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9082 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9083 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9084 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9085 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9086 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9087 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9088 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9089 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9090 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9091 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9092 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9093 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9094 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9095 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9096 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9097 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9098 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9099 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9100 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9101 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9102 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9103 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9104 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9105 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9106 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9107 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9108 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9109 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9110 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9111 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9112 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9113 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9114 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9115 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9116 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9117 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9118 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9119 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9120 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9121 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9122 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9123 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9124 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9125 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9126 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9127 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9128 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9129 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9130 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9131 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9132 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9133 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9134 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9135 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9136 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9137 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9138 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9139 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9140 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9141 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9142 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9143 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9144 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9145 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9146 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9147 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9148 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9149 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9150 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9151 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9152 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9153 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9154 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9155 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9156 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9157 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9158 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9159 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9160 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9161 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9162 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9163 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9164 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9165 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9166 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9167 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9168 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9169 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9170 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9171 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9172 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9173 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9174 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9175 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9176 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9177 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9178 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9179 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9180 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9181 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9182 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9183 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9184 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9185 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9186 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9187 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9188 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9189 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9190 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9191 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9192 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9193 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9194 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9195 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9196 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9197 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9198 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9199 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9200 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9201 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9202 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9203 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9204 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9205 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9206 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9207 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9208 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9209 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9210 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9211 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9212 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9213 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9214 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9215 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9216 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9217 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9218 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9219 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9220 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9221 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9222 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9223 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9224 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9225 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9226 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9227 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9228 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9229 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9230 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9231 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9232 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9233 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9234 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9235 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9236 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9237 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9238 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9239 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9240 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9241 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9242 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9243 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9244 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9245 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9246 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9247 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9248 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9249 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9250 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9251 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9252 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9253 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9254 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9255 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9256 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9257 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9258 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9259 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9260 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9261 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9262 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9263 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9264 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9265 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9266 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9267 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9268 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9269 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9270 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9271 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9272 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9273 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9274 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9275 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9276 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9277 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9278 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9279 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9280 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9281 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9282 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9283 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9284 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9285 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9286 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9287 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9288 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9289 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9290 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9291 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9292 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9293 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9294 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9295 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9296 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9297 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9298 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9299 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9300 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9301 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9302 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9303 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9304 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9305 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9306 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9307 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9308 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9309 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9310 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9311 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9312 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9313 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9314 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9315 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9316 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9317 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9318 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9319 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9320 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9321 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9322 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9323 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9324 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9325 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9326 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9327 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9328 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9329 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9330 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9331 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9332 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9333 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9334 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9335 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9336 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9337 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9338 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9339 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9340 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9341 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9342 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9343 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9344 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9345 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9346 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9347 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9348 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9349 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9350 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9351 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9352 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9353 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9354 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9355 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9356 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9357 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9358 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9359 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9360 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9361 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9362 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9363 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9364 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9365 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9366 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9367 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9368 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9369 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9370 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9371 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9372 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9373 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9374 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9375 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9376 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9377 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9378 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9379 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9380 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9381 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9382 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9383 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9384 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9385 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9386 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9387 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9388 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9389 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9390 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9391 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9392 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9393 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9394 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9395 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9396 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9397 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9398 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9399 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9400 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9401 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9402 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9403 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9404 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9405 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9406 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9407 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9408 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9409 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9410 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9411 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9412 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9413 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9414 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9415 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9416 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9417 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9418 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9419 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9420 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9421 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9422 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9423 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9424 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9425 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9426 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9427 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9428 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9429 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9430 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9431 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9432 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9433 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9434 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9435 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9436 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9437 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9438 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9439 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9440 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9441 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9442 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9443 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9444 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9445 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9446 10bitdac_layout_0/inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9447 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 10bitdac_layout_0/inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9448 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9449 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9450 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9451 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9452 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9453 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9454 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9455 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9456 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9457 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9458 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9459 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 10bitdac_layout_0/inp2 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9460 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9461 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9462 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9463 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_vref5 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
C0 10bitdac_layout_0/d5 10bitdac_layout_0/d3 29.02fF
C1 10bitdac_layout_0/d3 10bitdac_layout_0/9bitdac_layout_1/d2 67.70fF
C2 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 12.72fF
C3 10bitdac_layout_0/d4 10bitdac_layout_0/d3 129.84fF
C4 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 12.72fF
C5 10bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 5.86fF
C6 10bitdac_layout_0/9bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 3.29fF
C7 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/x2_vref1 19.77fF
C8 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 2.44fF
C9 10bitdac_layout_0/d6 10bitdac_layout_0/d7 23.66fF
C10 10bitdac_layout_0/9bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_vref1 3.09fF
C11 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 2.44fF
C12 10bitdac_layout_0/d0 vdd 53.48fF
C13 10bitdac_layout_0/d1 vdd 42.81fF
C14 10bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 8.21fF
C15 10bitdac_layout_0/d0 10bitdac_layout_0/d5 11.54fF
C16 10bitdac_layout_0/d2 vdd 8.89fF
C17 10bitdac_layout_0/d5 10bitdac_layout_0/d1 5.05fF
C18 10bitdac_layout_0/d0 10bitdac_layout_0/9bitdac_layout_1/d2 16.85fF
C19 10bitdac_layout_0/d4 10bitdac_layout_0/d0 5.09fF
C20 10bitdac_layout_0/d1 10bitdac_layout_0/9bitdac_layout_1/d2 49.96fF
C21 10bitdac_layout_0/d4 10bitdac_layout_0/d1 7.44fF
C22 10bitdac_layout_0/d0 10bitdac_layout_0/d3 6.80fF
C23 10bitdac_layout_0/d2 10bitdac_layout_0/d5 3.34fF
C24 10bitdac_layout_0/d1 10bitdac_layout_0/d3 36.27fF
C25 10bitdac_layout_0/d4 10bitdac_layout_0/d2 20.08fF
C26 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_out_v 2.44fF
C27 10bitdac_layout_0/d2 10bitdac_layout_0/d3 67.70fF
C28 10bitdac_layout_0/d5 10bitdac_layout_0/d7 4.02fF
C29 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 3.09fF
C30 10bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 3.14fF
C31 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x2_vref1 12.72fF
C32 10bitdac_layout_0/d5 10bitdac_layout_0/d6 56.74fF
C33 10bitdac_layout_0/d4 10bitdac_layout_0/d6 22.94fF
C34 10bitdac_layout_0/9bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 19.77fF
C35 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/x1_out_v 34.19fF
C36 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/x2_vref1 12.72fF
C37 10bitdac_layout_0/d0 10bitdac_layout_0/d1 179.55fF
C38 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/x1_out_v 34.19fF
C39 10bitdac_layout_0/d2 10bitdac_layout_0/d0 16.90fF
C40 10bitdac_layout_0/d2 10bitdac_layout_0/d1 49.96fF
C41 vdd 10bitdac_layout_0/9bitdac_layout_1/d2 8.96fF
C42 10bitdac_layout_0/9bitdac_layout_0/x2_vref1 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/x1_out_v 3.29fF
C43 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/x1_out_v 2.44fF
C44 10bitdac_layout_0/d3 vdd 6.90fF
C45 10bitdac_layout_0/d5 10bitdac_layout_0/9bitdac_layout_1/d2 3.34fF
C46 10bitdac_layout_0/d4 10bitdac_layout_0/d5 95.86fF
C47 10bitdac_layout_0/d4 10bitdac_layout_0/9bitdac_layout_1/d2 20.08fF
C48 10bitdac_layout_0/d0 10bitdac_layout_0/d6 28.63fF
C49 10bitdac_layout_0/d1 10bitdac_layout_0/d6 15.27fF
C50 vdd 0 1922.01fF
C51 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C52 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C53 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C54 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C55 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 2.08fF
C56 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C57 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C58 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C59 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C60 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C61 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C62 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C63 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C64 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 2.08fF
C65 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C66 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C67 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C68 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C69 10bitdac_layout_0/9bitdac_layout_1/x1_vref5 0 2.19fF
C70 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C71 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C72 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C73 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C74 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 2.08fF
C75 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C76 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C77 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C78 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C79 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C80 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C81 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C82 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C83 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 2.08fF
C84 10bitdac_layout_0/d0 0 858.43fF
C85 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C86 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C87 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C88 10bitdac_layout_0/9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C89 10bitdac_layout_0/d5 0 506.12fF
C90 10bitdac_layout_0/d6 0 310.51fF
C91 10bitdac_layout_0/d7 0 169.86fF
C92 10bitdac_layout_0/x1_vref5 0 2.09fF
C93 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C94 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C95 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C96 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C97 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 2.08fF
C98 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C99 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C100 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C101 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C102 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C103 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C104 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C105 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C106 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 2.08fF
C107 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C108 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C109 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C110 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C111 10bitdac_layout_0/9bitdac_layout_0/x1_vref5 0 2.19fF
C112 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C113 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C114 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C115 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C116 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 2.08fF
C117 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C118 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C119 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C120 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C121 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C122 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C123 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C124 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C125 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 2.08fF
C126 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C127 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C128 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C129 10bitdac_layout_0/9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C130 m1_104169_26312# 0 1129.51fF **FLOATING

V1 vdd 0 dc 3.3V
V2 d0 0 PULSE 0 1.8 0ns 1p 1p 5u 10u
V3 d1 0 PULSE 0 1.8 0ns 1p 1p 10u 20u
V4 inp2 0 dc 0V
V5 inp1 0 dc 3.3V
V6 d2 0 PULSE 0 1.8 0ns 1p 1p 20u 40u
V7 d3 0 PULSE 0 1.8 0ns 1p 1p 40u 80u
V8 d4 0 PULSE 0 1.8 0ns 1p 1p 80u 160u
V9 d5 0 PULSE 0 1.8 0ns 1p 1p 160u 320u
V10 d6 0 PULSE 0 1.8 0 1p 1p 320u 640u
V11 d7 0 PULSE 0 1.8 0 1p 1p 640u 1280u
V12 d8 0 PULSE 0 1.8 0 1p 1p 1280u 2560u
V13 d9 0 PULSE 0 1.8 0 1p 1p 2560u 5120u

.tran 2u 5120u
.control
run 
plot d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 out_v
plot out_v
.endc
.end
