magic
tech sky130A
timestamp 1625518311
<< metal1 >>
rect -984 12417 -496 12449
rect -984 11818 12410 12417
rect -984 -1163 12375 11818
rect -984 -1226 -464 -1163
rect 11855 -1226 12375 -1163
<< metal3 >>
rect -984 12417 -496 12449
rect -984 11818 12410 12417
rect -984 11706 12375 11818
rect -984 -442 -260 11706
rect 11803 -442 12375 11706
rect -984 -1163 12375 -442
rect -984 -1226 -464 -1163
rect 11855 -1226 12375 -1163
<< end >>
