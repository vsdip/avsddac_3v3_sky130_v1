* SPICE3 file created from res500_layout.ext - technology: sky130A
* Resistor value test

* Include SkyWater sky130 device models
.lib "../sky130_fd_pr/models/sky130.lib.spice" tt


* Simple voltage across a modeled device resistor
V1 0 A DC 1.8

X0 0 A 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24


.control
op lin 0 3.3
run
echo resistance
print V(A)/V1#branch
quit
.endc
.end
