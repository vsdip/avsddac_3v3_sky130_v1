magic
tech sky130A
timestamp 1616473885
<< locali >>
rect 200 654 1127 655
rect 1315 654 1507 655
rect 200 635 1507 654
rect 200 634 1436 635
rect 200 533 221 634
rect 1126 633 1316 634
rect 85 369 110 493
rect 200 432 220 533
rect 1489 530 1507 635
rect 75 219 100 269
rect 201 219 220 432
rect 1712 427 1734 428
rect 1712 408 3080 427
rect 1712 395 1734 408
rect 1566 390 1734 395
rect 1566 371 1572 390
rect 1590 371 1734 390
rect 1566 365 1734 371
rect 1566 364 1732 365
rect 389 329 408 331
rect 75 199 220 219
rect 384 205 408 329
rect 3055 288 3080 408
rect 75 145 100 199
rect 336 86 364 92
rect 336 85 340 86
rect 195 66 340 85
rect 359 66 364 86
rect 384 84 409 205
rect 454 88 482 91
rect 1499 88 1528 153
rect 3136 148 3251 153
rect 3136 129 3140 148
rect 3158 129 3251 148
rect 3136 121 3251 129
rect 454 87 1528 88
rect 195 65 364 66
rect 74 0 102 46
rect 195 0 218 65
rect 336 59 364 65
rect 386 64 409 84
rect 452 84 1528 87
rect 452 64 458 84
rect 477 64 1528 84
rect 386 62 408 64
rect 334 4 361 10
rect 334 2 338 4
rect 74 -21 218 0
rect 273 -15 338 2
rect 357 -15 361 4
rect 273 -20 361 -15
rect 74 -170 102 -21
rect 273 -101 295 -20
rect 334 -23 361 -20
rect 385 6 408 62
rect 454 63 1528 64
rect 454 62 1524 63
rect 454 58 482 62
rect 1916 39 2031 90
rect 447 6 476 11
rect 385 -13 409 6
rect 447 5 1522 6
rect 385 -60 408 -13
rect 447 -14 451 5
rect 470 -12 1522 5
rect 470 -14 476 -12
rect 931 -13 1294 -12
rect 447 -22 476 -14
rect 348 -82 408 -60
rect 96 -171 102 -170
rect 83 -316 130 -271
rect 100 -356 130 -316
rect 272 -354 295 -101
rect 384 -353 408 -82
rect 1502 -111 1522 -12
rect 3078 -241 3098 -86
rect 2322 -243 2441 -242
rect 2540 -243 2659 -242
rect 2762 -243 2881 -242
rect 2980 -243 3099 -241
rect 2101 -244 3099 -243
rect 1762 -246 1881 -245
rect 1990 -246 3099 -244
rect 1578 -254 3099 -246
rect 1578 -272 1585 -254
rect 1602 -269 3099 -254
rect 1602 -270 2994 -269
rect 1602 -271 2331 -270
rect 2432 -271 2551 -270
rect 2647 -271 2766 -270
rect 2875 -271 2994 -270
rect 1602 -272 2109 -271
rect 1578 -273 1995 -272
rect 1578 -274 1767 -273
rect 1876 -274 1995 -273
rect 1578 -275 1650 -274
rect 179 -356 295 -354
rect 388 -356 408 -353
rect 100 -374 295 -356
rect 100 -375 165 -374
rect 100 -454 130 -375
rect -5 -570 20 -493
rect 792 -549 976 -548
rect 1517 -549 1534 -486
rect 166 -550 190 -549
rect 274 -550 1534 -549
rect 166 -566 1534 -550
rect 166 -567 1317 -566
rect 165 -568 797 -567
rect 952 -568 1317 -567
rect 165 -569 352 -568
rect 165 -570 190 -569
rect -5 -587 190 -570
rect -5 -617 20 -587
<< viali >>
rect 1572 371 1590 390
rect 340 66 359 86
rect 3140 129 3158 148
rect 458 64 477 84
rect 338 -15 357 4
rect 451 -14 470 5
rect 1585 -272 1602 -254
<< metal1 >>
rect 801 563 811 600
rect 801 562 841 563
rect 801 557 847 562
rect 801 523 814 557
rect 842 523 847 557
rect 801 518 847 523
rect 2371 317 2432 321
rect 2371 277 2389 317
rect 2426 277 2432 317
rect 2371 274 2432 277
rect 453 165 483 187
rect 453 136 454 165
rect 481 136 483 165
rect 453 115 483 136
rect 336 86 364 92
rect 454 88 482 91
rect 336 84 340 86
rect 335 66 340 84
rect 359 84 364 86
rect 452 84 483 88
rect 359 66 458 84
rect 335 64 458 66
rect 477 65 483 84
rect 477 64 482 65
rect 336 59 364 64
rect 454 58 482 64
rect 334 6 361 10
rect 447 6 476 11
rect 334 5 476 6
rect 334 4 451 5
rect 334 -15 338 4
rect 357 -13 451 4
rect 357 -15 361 -13
rect 334 -23 361 -15
rect 447 -14 451 -13
rect 470 -14 476 5
rect 447 -22 476 -14
rect 822 -84 866 -77
rect 822 -119 831 -84
rect 860 -119 866 -84
rect 822 -124 866 -119
rect 2015 -86 2056 -54
rect 2015 -113 2019 -86
rect 2046 -113 2056 -86
rect 2015 -125 2056 -113
rect 2029 -126 2056 -125
rect 471 -476 501 -452
rect 498 -505 501 -476
rect 471 -524 501 -505
<< via1 >>
rect 814 523 842 557
rect 2389 277 2426 317
rect 454 136 481 165
rect 831 -119 860 -84
rect 2019 -113 2046 -86
rect 471 -505 498 -476
<< metal2 >>
rect 811 606 853 617
rect 811 568 815 606
rect 848 568 853 606
rect 811 565 853 568
rect 811 557 847 565
rect 811 523 814 557
rect 842 523 847 557
rect 811 517 847 523
rect 2383 369 2433 376
rect 2383 324 2390 369
rect 2426 324 2433 369
rect 2383 317 2433 324
rect 2383 277 2389 317
rect 2426 277 2433 317
rect 2383 274 2433 277
rect 436 165 484 169
rect 436 136 454 165
rect 481 136 484 165
rect 436 129 484 136
rect 436 -468 455 129
rect 828 -38 866 -33
rect 828 -73 832 -38
rect 861 -73 866 -38
rect 828 -84 866 -73
rect 2000 -81 2021 -80
rect 828 -119 831 -84
rect 860 -119 866 -84
rect 1955 -85 2047 -81
rect 828 -124 866 -119
rect 1950 -86 2047 -85
rect 1950 -113 2019 -86
rect 2046 -89 2047 -86
rect 2046 -113 2048 -89
rect 1950 -116 2048 -113
rect 1950 -119 2047 -116
rect 1950 -342 1974 -119
rect 2000 -120 2021 -119
rect 1950 -457 1975 -342
rect 436 -471 461 -468
rect 436 -476 501 -471
rect 436 -505 471 -476
rect 498 -505 501 -476
rect 436 -511 501 -505
rect 437 -625 461 -511
rect 1951 -625 1975 -457
rect 437 -642 1975 -625
rect 437 -649 1948 -642
<< via2 >>
rect 815 568 848 606
rect 2390 324 2426 369
rect 832 -73 861 -38
<< metal3 >>
rect 810 708 864 713
rect 810 662 815 708
rect 853 662 864 708
rect 810 658 864 662
rect 811 617 851 658
rect 811 606 853 617
rect 811 568 815 606
rect 848 568 853 606
rect 811 565 853 568
rect 811 563 847 565
rect 2383 474 2434 478
rect 2383 434 2391 474
rect 2425 434 2434 474
rect 2383 429 2434 434
rect 2383 369 2433 429
rect 2383 324 2390 369
rect 2426 324 2433 369
rect 2383 321 2433 324
rect 828 45 873 52
rect 828 12 833 45
rect 867 12 873 45
rect 828 9 873 12
rect 828 -38 872 9
rect 828 -73 832 -38
rect 861 -73 872 -38
rect 828 -77 872 -73
<< via3 >>
rect 815 662 853 708
rect 2391 434 2425 474
rect 833 12 867 45
<< metal4 >>
rect 1094 713 2021 714
rect 2244 713 2435 715
rect 811 708 2435 713
rect 811 662 815 708
rect 853 662 2435 708
rect 811 661 2435 662
rect 811 660 2252 661
rect 811 659 1095 660
rect 2016 659 2252 660
rect 872 51 927 659
rect 2383 478 2432 661
rect 2383 474 2434 478
rect 2383 434 2391 474
rect 2425 434 2434 474
rect 2383 429 2434 434
rect 828 45 927 51
rect 828 12 833 45
rect 867 12 927 45
rect 828 11 927 12
rect 828 9 886 11
use res500_layout  res500_layout_0
timestamp 1615766096
transform 0 1 144 -1 0 299
box 109 -144 299 -45
use res500_layout  res500_layout_1
timestamp 1615766096
transform 0 1 144 -1 0 -17
box 109 -144 299 -45
use res500_layout  res500_layout_2
timestamp 1615766096
transform 0 1 148 -1 0 523
box 109 -144 299 -45
use res250_layout  res250_layout_0
timestamp 1615764517
transform 0 1 170 -1 0 -299
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 366 0 1 25
box 20 86 1230 590
use switch_layout  switch_layout_1
timestamp 1615739263
transform 1 0 382 0 1 -615
box 20 86 1230 590
use switch_layout  switch_layout_2
timestamp 1615739263
transform 1 0 1934 0 1 -217
box 20 86 1230 590
<< labels >>
rlabel locali 100 408 100 408 1 vref1
rlabel locali 98 206 98 206 1 x1_inp1
rlabel locali 80 -64 80 -64 1 x1_inp2
rlabel locali 122 -365 122 -365 1 x2_inp1
rlabel locali 3 -577 3 -577 1 vref5
rlabel locali 390 -81 390 -81 1 d0
rlabel locali 1934 60 1934 60 1 d1
rlabel locali 1651 377 1651 377 1 x1_vout
rlabel locali 1765 -260 1765 -260 1 x2_vout
rlabel locali 3198 137 3198 137 1 out_v
rlabel metal4 1118 687 1118 687 1 vdd!
rlabel metal2 1031 -637 1031 -637 1 gnd!
<< end >>
