magic
tech sky130A
timestamp 1616493856
<< locali >>
rect 22885 25777 45390 25781
rect 47680 25777 48092 25779
rect 22885 25760 48092 25777
rect 22885 25686 22912 25760
rect 47682 25758 48092 25760
rect 22885 25667 22888 25686
rect 22906 25667 22912 25686
rect 22885 25663 22912 25667
rect 48074 25733 48092 25758
rect 10595 25639 10873 25640
rect 10595 25637 18730 25639
rect 10185 25636 18730 25637
rect 10185 25629 24077 25636
rect 10185 25615 10196 25629
rect 10186 25609 10196 25615
rect 10220 25617 24077 25629
rect 10220 25615 10695 25617
rect 10220 25609 10226 25615
rect 10186 25605 10226 25609
rect 22884 25596 22909 25598
rect 22884 25577 22888 25596
rect 22906 25577 22909 25596
rect 398 25313 427 25336
rect 398 25295 405 25313
rect 423 25295 427 25313
rect 398 25293 427 25295
rect 10191 25207 10228 25216
rect 10191 25187 10196 25207
rect 10220 25187 10228 25207
rect 10191 24780 10228 25187
rect 22884 24908 22909 25577
rect 24049 25331 24077 25617
rect 24046 25324 24079 25331
rect 24046 25302 24053 25324
rect 24075 25302 24079 25324
rect 24046 25297 24079 25302
rect 24049 25295 24077 25297
rect 10190 13096 10230 24780
rect 22884 13737 22908 24908
rect 48074 24601 48095 25733
rect 48073 13811 48095 24601
rect 48073 13790 48098 13811
rect 21561 13366 21581 13702
rect 21561 13348 21562 13366
rect 21579 13348 21581 13366
rect 21561 13341 21581 13348
rect 45188 13382 45234 13696
rect 45188 13356 45197 13382
rect 45221 13356 45234 13382
rect 45188 13329 45234 13356
rect 21555 13259 21582 13263
rect 21555 13241 21560 13259
rect 21577 13241 21582 13259
rect 21555 13236 21582 13241
rect 10190 13081 10233 13096
rect 10193 1405 10233 13081
rect 21558 12703 21582 13236
rect 21555 12193 21582 12703
rect 21551 11964 21582 12193
rect 45188 13205 45217 13230
rect 45188 13179 45191 13205
rect 45215 13179 45217 13205
rect 10193 1156 10236 1405
rect 10191 1144 10236 1156
rect 10191 940 10234 1144
rect 10300 1092 10351 1179
rect 10388 940 10439 987
rect 10191 895 10442 940
rect 10193 894 10442 895
rect 10646 -585 10676 24
rect 12185 -513 12215 96
rect 13855 -409 13885 220
rect 15552 -318 15582 367
rect 17173 -221 17203 510
rect 18904 -150 18934 728
rect 21551 646 21577 11964
rect 33984 1130 34013 1177
rect 21546 -54 21579 646
rect 24251 22 24286 27
rect 39271 25 39319 331
rect 40845 26 40894 501
rect 42560 216 42591 699
rect 42560 49 42595 216
rect 42560 43 42601 49
rect 42560 36 42566 43
rect 24251 0 24260 22
rect 24280 0 24286 22
rect 24251 -5 24286 0
rect 39270 18 39320 25
rect 39270 -12 39277 18
rect 39310 -12 39320 18
rect 40844 19 40895 26
rect 40844 4 40851 19
rect 39270 -19 39320 -12
rect 39271 -22 39319 -19
rect 40845 -20 40851 4
rect 40888 4 40895 19
rect 42563 10 42566 36
rect 42593 10 42601 43
rect 42563 4 42601 10
rect 40888 -20 40894 4
rect 42563 -2 42595 4
rect 40845 -24 40894 -20
rect 44146 -51 44821 -49
rect 45188 -51 45217 13179
rect 46516 13048 46556 13767
rect 48075 13661 48098 13790
rect 48160 13521 48260 13526
rect 48160 13498 48164 13521
rect 48184 13498 48260 13521
rect 48160 13494 48260 13498
rect 46965 13415 46990 13461
rect 48086 13182 48107 13285
rect 48086 13060 48109 13182
rect 48086 13050 48106 13060
rect 46770 13048 48106 13050
rect 46516 13015 48106 13048
rect 46516 13013 46781 13015
rect 44146 -54 45217 -51
rect 21545 -84 45217 -54
rect 21545 -86 42555 -84
rect 42613 -86 45217 -84
rect 21545 -93 21618 -86
rect 44146 -92 45217 -86
rect 42560 -124 42591 -119
rect 18900 -152 31660 -150
rect 42560 -152 42562 -124
rect 18900 -157 42562 -152
rect 42589 -136 42591 -124
rect 42589 -157 42597 -136
rect 18900 -181 42597 -157
rect 18900 -183 42589 -181
rect 18900 -186 31660 -183
rect 18904 -190 18934 -186
rect 17175 -234 17203 -221
rect 40844 -220 40895 -210
rect 40844 -230 40852 -220
rect 22140 -232 40852 -230
rect 19650 -234 40852 -232
rect 17175 -259 40852 -234
rect 40889 -232 40895 -220
rect 40889 -259 40894 -232
rect 17175 -260 40894 -259
rect 17175 -262 40879 -260
rect 17175 -264 35395 -262
rect 17175 -266 22152 -264
rect 17175 -267 19671 -266
rect 17224 -268 19671 -267
rect 15549 -322 18342 -318
rect 21082 -322 28711 -320
rect 15549 -324 32526 -322
rect 15549 -330 36347 -324
rect 39271 -330 39319 -326
rect 15549 -331 39319 -330
rect 15549 -348 39279 -331
rect 15552 -352 15582 -348
rect 18323 -352 39279 -348
rect 21082 -356 39279 -352
rect 28683 -358 39279 -356
rect 32504 -360 39279 -358
rect 39267 -361 39279 -360
rect 39312 -361 39319 -331
rect 39267 -365 39319 -361
rect 13849 -411 16864 -409
rect 13849 -417 37682 -411
rect 13849 -435 37653 -417
rect 37675 -433 37682 -417
rect 37675 -435 37681 -433
rect 13849 -438 37681 -435
rect 13855 -443 13885 -438
rect 37645 -442 37681 -438
rect 35897 -513 35931 -511
rect 12185 -514 35931 -513
rect 12185 -531 35904 -514
rect 35925 -531 35931 -514
rect 12185 -534 29313 -531
rect 12185 -535 19795 -534
rect 35897 -536 35931 -531
rect 23498 -585 24287 -580
rect 10643 -586 13876 -585
rect 20313 -586 24287 -585
rect 10643 -587 24287 -586
rect 10643 -607 24259 -587
rect 24279 -607 24287 -587
rect 10643 -612 24287 -607
rect 10643 -615 23546 -612
rect 10712 -616 13225 -615
rect 13867 -616 20325 -615
<< viali >>
rect 22888 25667 22906 25686
rect 10196 25609 10220 25629
rect 22888 25577 22906 25596
rect 405 25295 423 25313
rect 404 25208 422 25226
rect 10196 25187 10220 25207
rect 24053 25302 24075 25324
rect 24057 25201 24079 25223
rect 21562 13348 21579 13366
rect 45197 13356 45221 13382
rect 21560 13241 21577 13259
rect 45191 13179 45215 13205
rect 24260 0 24280 22
rect 39277 -12 39310 18
rect 40851 -20 40888 19
rect 42566 10 42593 43
rect 48164 13498 48184 13521
rect 42562 -157 42589 -124
rect 40852 -259 40889 -220
rect 39279 -361 39312 -331
rect 37653 -435 37675 -417
rect 35904 -531 35925 -514
rect 24259 -607 24279 -587
<< metal1 >>
rect 22883 25686 22912 25692
rect 22882 25667 22888 25686
rect 22906 25667 22912 25686
rect 22882 25663 22912 25667
rect 10188 25629 10225 25638
rect 10188 25609 10196 25629
rect 10220 25609 10225 25629
rect 398 25313 427 25328
rect 398 25295 405 25313
rect 423 25295 427 25313
rect 398 25226 427 25295
rect 398 25208 404 25226
rect 422 25208 427 25226
rect 398 25202 427 25208
rect 10188 25207 10225 25609
rect 22884 25596 22911 25663
rect 22883 25577 22888 25596
rect 22906 25577 22911 25596
rect 22883 25570 22911 25577
rect 24046 25329 24079 25331
rect 24046 25324 24084 25329
rect 24046 25302 24053 25324
rect 24075 25302 24084 25324
rect 24046 25297 24084 25302
rect 24050 25228 24084 25297
rect 10188 25187 10196 25207
rect 10220 25187 10225 25207
rect 24049 25223 24084 25228
rect 24049 25201 24057 25223
rect 24079 25206 24084 25223
rect 24079 25201 24082 25206
rect 24049 25194 24082 25201
rect 10188 25179 10225 25187
rect 47396 13677 47440 13683
rect 47396 13651 47412 13677
rect 47439 13651 47440 13677
rect 47396 13645 47440 13651
rect 48160 13521 48193 13526
rect 48160 13498 48164 13521
rect 48184 13498 48193 13521
rect 48160 13493 48193 13498
rect 45181 13382 45234 13396
rect 21558 13371 21581 13379
rect 21558 13366 21582 13371
rect 21558 13348 21562 13366
rect 21579 13348 21582 13366
rect 21558 13343 21582 13348
rect 45181 13356 45197 13382
rect 45221 13356 45234 13382
rect 21558 13263 21581 13343
rect 21555 13259 21581 13263
rect 21555 13241 21560 13259
rect 21577 13241 21581 13259
rect 21555 13236 21581 13241
rect 21558 13235 21581 13236
rect 45181 13205 45234 13356
rect 47024 13290 47080 13315
rect 47024 13262 47035 13290
rect 47064 13262 47080 13290
rect 47024 13246 47080 13262
rect 45181 13179 45191 13205
rect 45215 13179 45234 13205
rect 45181 13170 45234 13179
rect 24251 23 24286 27
rect 24251 22 24287 23
rect 24251 0 24260 22
rect 24280 0 24287 22
rect 24251 -5 24287 0
rect 24256 -581 24287 -5
rect 35899 -511 35929 86
rect 37644 -390 37682 218
rect 42561 49 42593 63
rect 42561 43 42601 49
rect 39270 18 39320 25
rect 39270 -12 39277 18
rect 39310 -12 39320 18
rect 40844 21 40895 26
rect 40844 19 40896 21
rect 40844 4 40851 19
rect 39270 -19 39320 -12
rect 39271 -331 39319 -19
rect 40847 -20 40851 4
rect 40888 -20 40896 19
rect 40847 -220 40896 -20
rect 42561 10 42566 43
rect 42593 10 42601 43
rect 42561 4 42601 10
rect 42561 -103 42593 4
rect 42557 -124 42593 -103
rect 42557 -157 42562 -124
rect 42589 -136 42593 -124
rect 42589 -157 42597 -136
rect 42557 -181 42597 -157
rect 42557 -189 42589 -181
rect 40847 -259 40852 -220
rect 40889 -259 40896 -220
rect 40847 -267 40896 -259
rect 39271 -346 39279 -331
rect 39270 -361 39279 -346
rect 39312 -361 39319 -331
rect 39270 -365 39319 -361
rect 37644 -411 37680 -390
rect 37644 -417 37682 -411
rect 37644 -435 37653 -417
rect 37675 -433 37682 -417
rect 37675 -435 37681 -433
rect 37644 -436 37681 -435
rect 37645 -442 37681 -436
rect 35897 -514 35931 -511
rect 35897 -531 35904 -514
rect 35925 -531 35931 -514
rect 35897 -536 35931 -531
rect 24253 -587 24287 -581
rect 24253 -607 24259 -587
rect 24279 -607 24287 -587
rect 24253 -612 24287 -607
<< via1 >>
rect 47412 13651 47439 13677
rect 47035 13262 47064 13290
<< metal2 >>
rect 12145 25455 12576 25460
rect 12145 25453 29141 25455
rect 12145 25427 29200 25453
rect 12145 25425 29141 25427
rect 12560 25424 29141 25425
rect 47405 13718 47440 13723
rect 47405 13690 47408 13718
rect 47436 13690 47440 13718
rect 47405 13677 47440 13690
rect 47405 13651 47412 13677
rect 47439 13651 47440 13677
rect 47405 13646 47440 13651
rect 46967 13293 47073 13296
rect 46957 13290 47073 13293
rect 46957 13262 47035 13290
rect 47064 13262 47073 13290
rect 46957 13250 47073 13262
rect 46957 13120 46977 13250
rect 45506 13119 46979 13120
rect 45250 13101 46979 13119
rect 45250 13100 46015 13101
rect 45250 13099 45507 13100
<< via2 >>
rect 47408 13690 47436 13718
<< metal3 >>
rect 47405 13765 47445 13769
rect 47405 13733 47410 13765
rect 47442 13733 47445 13765
rect 47405 13728 47445 13733
rect 47405 13718 47440 13728
rect 47405 13690 47408 13718
rect 47436 13690 47440 13718
rect 47405 13686 47440 13690
<< via3 >>
rect 47410 13733 47442 13765
<< metal4 >>
rect 11881 25748 24882 25750
rect 11376 25717 24882 25748
rect 11376 25716 11904 25717
rect 11382 25311 11424 25716
rect 24846 25157 24881 25717
rect 45667 14035 47445 14070
rect 47408 13795 47445 14035
rect 47405 13792 47445 13795
rect 47405 13765 47444 13792
rect 47405 13733 47410 13765
rect 47442 13733 47444 13765
rect 47405 13730 47444 13733
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 10196 0 1 1151
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 46957 0 1 13155
box 20 86 1230 590
use 7bitdac_layout  7bitdac_layout_1
timestamp 1616488517
transform 1 0 23779 0 1 1222
box -126 -1228 22781 24343
use 7bitdac_layout  7bitdac_layout_0
timestamp 1616488517
transform 1 0 126 0 1 1228
box -126 -1228 22781 24343
<< labels >>
rlabel locali 10326 1132 10326 1132 1 x1_vref5
rlabel locali 10406 934 10406 934 1 x2_vref1
rlabel locali 402 25332 402 25332 1 inp1
rlabel locali 33997 1147 33997 1147 1 inp2
rlabel locali 46976 13431 46976 13431 1 d7
rlabel locali 48226 13507 48226 13507 1 out_v
rlabel locali 48088 13772 48088 13772 1 x1_out_v
rlabel locali 48100 13194 48100 13194 1 x2_out_v
rlabel metal2 46989 13270 46989 13270 1 gnd!
rlabel metal4 47432 13777 47432 13777 1 vdd!
rlabel locali 21563 22 21563 22 1 d6
rlabel locali 18921 -109 18921 -109 1 d5
rlabel locali 17182 306 17182 306 1 d4
rlabel locali 15566 243 15566 243 1 d3
rlabel locali 13868 76 13868 76 1 d2
rlabel locali 12198 20 12198 20 1 d1
rlabel locali 10658 -32 10658 -32 1 d0
<< end >>
