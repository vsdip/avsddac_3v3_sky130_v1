magic
tech sky130A
magscale 1 2
timestamp 1624221218
<< checkpaint >>
rect -1688 -58952 206316 56030
<< locali >>
rect 796 53914 852 54034
rect 198700 29356 204742 29418
rect 195658 29180 196142 29254
rect 195658 28902 195742 29180
rect 195658 28868 195685 28902
rect 195719 28868 195742 28902
rect 195658 28848 195742 28868
rect 195664 28608 195734 28638
rect 195664 28574 195683 28608
rect 195717 28574 195734 28608
rect 195664 22018 195734 28574
rect 204674 24878 204742 29356
rect 204672 24802 204742 24878
rect 195664 21966 195744 22018
rect 165972 5160 166028 5278
rect 166150 4802 166236 4972
rect 166150 4768 166180 4802
rect 166214 4768 166236 4802
rect 166150 4766 166236 4768
rect 169778 2000 169812 2036
rect 169778 1990 169826 2000
rect 166148 1950 166242 1962
rect 166148 1928 166176 1950
rect 166146 1916 166176 1928
rect 166210 1916 166242 1950
rect 166146 1896 166242 1916
rect 166146 1212 166230 1896
rect 166138 1199 166230 1212
rect 169778 1206 169812 1990
rect 173138 1268 173228 2234
rect 173138 1234 173160 1268
rect 173194 1234 173228 1268
rect 166138 1165 166150 1199
rect 166184 1165 166230 1199
rect 166138 1162 166230 1165
rect 166140 1160 166230 1162
rect 169774 1194 169832 1206
rect 173138 1202 173228 1234
rect 176554 1241 176612 2398
rect 179390 2076 179450 2602
rect 179390 1988 179466 2076
rect 176554 1207 176569 1241
rect 176603 1207 176612 1241
rect 169774 1160 169786 1194
rect 169820 1160 169832 1194
rect 176554 1192 176612 1207
rect 179394 1224 179466 1988
rect 179394 1190 179418 1224
rect 179452 1190 179466 1224
rect 179394 1170 179466 1190
rect 182738 1232 182788 2766
rect 182738 1198 182748 1232
rect 182782 1198 182788 1232
rect 182738 1180 182788 1198
rect 187976 1238 188046 2962
rect 187976 1204 187997 1238
rect 188031 1204 188046 1238
rect 187976 1176 188046 1204
rect 166140 1158 166208 1160
rect 169774 1150 169832 1160
rect 166788 1014 166860 1022
rect 169770 1018 169828 1032
rect 191468 1028 191536 1124
rect 166554 996 166870 1014
rect 166138 976 166186 978
rect 166138 942 166146 976
rect 166180 942 166186 976
rect 166554 962 166809 996
rect 166843 962 166870 996
rect 169770 984 169781 1018
rect 169815 984 169828 1018
rect 169770 972 169828 984
rect 179402 1008 179474 1028
rect 179402 974 179422 1008
rect 179456 974 179474 1008
rect 166554 942 166870 962
rect 166138 924 166186 942
rect 166138 268 166180 924
rect 166558 570 166598 942
rect 166788 940 166860 942
rect 169776 906 169812 972
rect 176554 941 176620 968
rect 169616 866 169812 906
rect 169620 758 169676 866
rect 169776 862 169812 866
rect 173132 878 173216 932
rect 173132 844 173156 878
rect 173190 844 173216 878
rect 169620 712 169678 758
rect 166558 530 166602 570
rect 166122 222 166180 268
rect 368 -2678 116520 -2670
rect 166122 -2678 166170 222
rect 166562 -1918 166602 530
rect 169624 6 169678 712
rect 169624 -34 169680 6
rect 169626 -746 169680 -34
rect 169626 -786 169682 -746
rect 169628 -1456 169682 -786
rect 173132 -916 173216 844
rect 169626 -1538 169682 -1456
rect 173130 -1006 173216 -916
rect 176554 907 176569 941
rect 176603 907 176620 941
rect 166562 -1946 166610 -1918
rect 368 -2716 166170 -2678
rect 368 -2720 116520 -2716
rect 368 -3772 424 -2720
rect 166568 -2818 166610 -1946
rect 166558 -2848 166630 -2818
rect 166558 -2882 166573 -2848
rect 166607 -2882 166630 -2848
rect 166558 -2900 166630 -2882
rect 169626 -2870 169680 -1538
rect 173130 -2778 173208 -1006
rect 173130 -2812 173156 -2778
rect 173190 -2812 173208 -2778
rect 173130 -2840 173208 -2812
rect 176554 -2780 176620 907
rect 179402 208 179474 974
rect 187972 992 188042 1022
rect 179398 122 179474 208
rect 182740 948 182788 972
rect 182740 914 182748 948
rect 182782 914 182788 948
rect 179398 -810 179462 122
rect 176554 -2814 176569 -2780
rect 176603 -2814 176620 -2780
rect 176554 -2842 176620 -2814
rect 179394 -886 179462 -810
rect 179394 -2750 179458 -886
rect 179394 -2784 179412 -2750
rect 179446 -2784 179458 -2750
rect 179394 -2836 179458 -2784
rect 182740 -2812 182788 914
rect 182738 -2816 182788 -2812
rect 182738 -2850 182746 -2816
rect 182780 -2850 182788 -2816
rect 182738 -2864 182788 -2850
rect 169626 -2904 169637 -2870
rect 169671 -2904 169680 -2870
rect 182740 -2880 182788 -2864
rect 187972 958 187993 992
rect 188027 958 188042 992
rect 187972 -2850 188042 958
rect 169626 -2916 169680 -2904
rect 187972 -2884 187991 -2850
rect 188025 -2884 188042 -2850
rect 191462 -2815 191536 1028
rect 191462 -2849 191479 -2815
rect 191513 -2849 191536 -2815
rect 191462 -2874 191536 -2849
rect 195668 -2862 195744 21966
rect 204672 190 204740 24802
rect 204862 -96 205056 -74
rect 204862 -130 204872 -96
rect 204906 -130 205056 -96
rect 204862 -144 205056 -130
rect 202362 -308 202584 -212
rect 204698 -996 204766 -552
rect 187972 -2908 188042 -2884
rect 195668 -2896 195690 -2862
rect 195724 -2896 195744 -2862
rect 195668 -2926 195744 -2896
rect 204054 -1054 204766 -996
rect 204054 -1060 204754 -1054
rect 195662 -3104 195738 -3078
rect 195662 -3138 195686 -3104
rect 195720 -3138 195738 -3104
rect 191448 -3223 191518 -3202
rect 191448 -3257 191467 -3223
rect 191501 -3257 191518 -3223
rect 187970 -3608 188038 -3590
rect 169616 -3652 169692 -3632
rect 169616 -3686 169633 -3652
rect 169667 -3686 169692 -3652
rect 169616 -3702 169692 -3686
rect 173128 -3690 173208 -3626
rect 182744 -3650 182790 -3614
rect 166560 -4454 166606 -4452
rect 166550 -4460 166618 -4454
rect 166550 -4490 166567 -4460
rect 166552 -4494 166567 -4490
rect 166601 -4494 166618 -4460
rect 166552 -4506 166618 -4494
rect 166566 -5002 166600 -4506
rect 169620 -4736 169674 -3702
rect 173128 -3724 173158 -3690
rect 173192 -3724 173208 -3690
rect 169618 -4752 169678 -4736
rect 169618 -4786 169635 -4752
rect 169669 -4786 169678 -4752
rect 169618 -4794 169678 -4786
rect 169624 -4944 169684 -4942
rect 169622 -4955 169684 -4944
rect 169622 -4989 169636 -4955
rect 169670 -4989 169684 -4955
rect 166566 -5020 166602 -5002
rect 169622 -5006 169684 -4989
rect 166566 -5022 166604 -5020
rect 166566 -5036 166600 -5022
rect 169624 -5536 169678 -5006
rect 173128 -5284 173208 -3724
rect 176548 -3690 176614 -3666
rect 176548 -3724 176567 -3690
rect 176601 -3724 176614 -3690
rect 173134 -6614 173202 -5524
rect 176548 -6294 176614 -3724
rect 179398 -3712 179462 -3658
rect 179398 -3746 179412 -3712
rect 179446 -3746 179462 -3712
rect 179398 -4462 179462 -3746
rect 182744 -3684 182748 -3650
rect 182782 -3684 182790 -3650
rect 179398 -4752 179466 -4462
rect 179402 -5508 179466 -4752
rect 179402 -5556 179470 -5508
rect 176548 -6328 176563 -6294
rect 176597 -6328 176614 -6294
rect 176548 -6356 176614 -6328
rect 179406 -6536 179470 -5556
rect 179402 -6602 179470 -6536
rect 173134 -6616 173248 -6614
rect 173134 -6656 173202 -6616
rect 176554 -6763 176626 -6732
rect 176554 -6797 176572 -6763
rect 176606 -6797 176626 -6763
rect 176554 -9876 176626 -6797
rect 179402 -9612 179466 -6602
rect 182744 -6958 182790 -3684
rect 187970 -3642 187991 -3608
rect 188025 -3642 188038 -3608
rect 182744 -7010 182802 -6958
rect 179402 -9646 179418 -9612
rect 179452 -9646 179466 -9612
rect 179402 -9660 179466 -9646
rect 179400 -9844 179470 -9830
rect 179400 -9878 179420 -9844
rect 179454 -9878 179470 -9844
rect 179400 -9896 179470 -9878
rect 179402 -9956 179470 -9896
rect 179406 -11952 179470 -9956
rect 179402 -12004 179470 -11952
rect 179402 -15108 179466 -12004
rect 182748 -14804 182802 -7010
rect 182748 -14818 182810 -14804
rect 182748 -14852 182762 -14818
rect 182796 -14852 182810 -14818
rect 182748 -14862 182810 -14852
rect 182748 -15050 182798 -15048
rect 182742 -15062 182802 -15050
rect 182742 -15096 182752 -15062
rect 182786 -15096 182802 -15062
rect 182742 -15108 182802 -15096
rect 182748 -15822 182798 -15108
rect 182748 -23716 182802 -15822
rect 182748 -23774 182806 -23716
rect 182752 -27720 182806 -23774
rect 187970 -26430 188038 -3642
rect 187970 -27264 188048 -26430
rect 191448 -27726 191518 -3257
rect 195662 -28022 195738 -3138
rect 195664 -28404 195738 -28022
rect 204054 -28274 204108 -1060
rect 198296 -28336 204108 -28274
rect 204054 -28338 204108 -28336
rect 195664 -28406 195778 -28404
rect 195664 -28488 195738 -28406
rect 165560 -52582 165620 -52438
<< viali >>
rect 195685 28868 195719 28902
rect 195683 28574 195717 28608
rect 166180 4768 166214 4802
rect 166176 1916 166210 1950
rect 173160 1234 173194 1268
rect 166150 1165 166184 1199
rect 176569 1207 176603 1241
rect 169786 1160 169820 1194
rect 179418 1190 179452 1224
rect 182748 1198 182782 1232
rect 187997 1204 188031 1238
rect 166146 942 166180 976
rect 166809 962 166843 996
rect 169781 984 169815 1018
rect 179422 974 179456 1008
rect 173156 844 173190 878
rect 176569 907 176603 941
rect 166573 -2882 166607 -2848
rect 173156 -2812 173190 -2778
rect 182748 914 182782 948
rect 176569 -2814 176603 -2780
rect 179412 -2784 179446 -2750
rect 182746 -2850 182780 -2816
rect 169637 -2904 169671 -2870
rect 187993 958 188027 992
rect 187991 -2884 188025 -2850
rect 191479 -2849 191513 -2815
rect 204872 -130 204906 -96
rect 195690 -2896 195724 -2862
rect 195686 -3138 195720 -3104
rect 191467 -3257 191501 -3223
rect 169633 -3686 169667 -3652
rect 166567 -4494 166601 -4460
rect 173158 -3724 173192 -3690
rect 169635 -4786 169669 -4752
rect 169636 -4989 169670 -4955
rect 176567 -3724 176601 -3690
rect 179412 -3746 179446 -3712
rect 182748 -3684 182782 -3650
rect 176563 -6328 176597 -6294
rect 176572 -6797 176606 -6763
rect 187991 -3642 188025 -3608
rect 179418 -9646 179452 -9612
rect 179420 -9878 179454 -9844
rect 182762 -14852 182796 -14818
rect 182752 -15096 182786 -15062
<< metal1 >>
rect 195658 28902 195742 28922
rect 195658 28868 195685 28902
rect 195719 28868 195742 28902
rect 195658 28608 195742 28868
rect 195658 28574 195683 28608
rect 195717 28574 195742 28608
rect 195658 28548 195742 28574
rect 166150 4802 166238 4810
rect 166150 4768 166180 4802
rect 166214 4768 166238 4802
rect 166150 1950 166238 4768
rect 166150 1916 166176 1950
rect 166210 1916 166238 1950
rect 166150 1896 166238 1916
rect 166798 1954 166838 3114
rect 166798 1844 166844 1954
rect 166138 1208 166206 1212
rect 166138 1199 166208 1208
rect 166138 1165 166150 1199
rect 166184 1165 166208 1199
rect 166138 1162 166208 1165
rect 166140 1158 166208 1162
rect 166140 976 166186 1158
rect 166802 1022 166844 1844
rect 173132 1268 173222 1334
rect 173132 1234 173160 1268
rect 173194 1234 173222 1268
rect 169774 1194 169832 1206
rect 169774 1160 169786 1194
rect 169820 1160 169832 1194
rect 169774 1150 169832 1160
rect 169778 1032 169814 1150
rect 166138 942 166146 976
rect 166180 942 166186 976
rect 166138 924 166186 942
rect 166788 996 166860 1022
rect 166788 962 166809 996
rect 166843 962 166860 996
rect 169770 1018 169828 1032
rect 169770 984 169781 1018
rect 169815 984 169828 1018
rect 169770 972 169828 984
rect 166788 940 166860 962
rect 173132 878 173222 1234
rect 176548 1241 176620 1292
rect 176548 1207 176569 1241
rect 176603 1207 176620 1241
rect 176548 941 176620 1207
rect 179402 1224 179470 1244
rect 179402 1190 179418 1224
rect 179452 1190 179470 1224
rect 179402 1008 179470 1190
rect 179402 974 179422 1008
rect 179456 974 179470 1008
rect 179402 948 179470 974
rect 182738 1232 182788 1256
rect 182738 1198 182748 1232
rect 182782 1198 182788 1232
rect 182738 948 182788 1198
rect 176548 907 176569 941
rect 176603 907 176620 941
rect 176548 884 176620 907
rect 182738 914 182748 948
rect 182782 914 182788 948
rect 187976 1238 188046 1266
rect 187976 1204 187997 1238
rect 188031 1204 188046 1238
rect 187976 992 188046 1204
rect 187976 958 187993 992
rect 188027 958 188046 992
rect 187976 934 188046 958
rect 182738 898 182788 914
rect 173132 844 173156 878
rect 173190 844 173222 878
rect 173132 806 173222 844
rect 203326 230 203420 238
rect 203326 178 203361 230
rect 203413 178 203420 230
rect 203326 164 203420 178
rect 204864 -96 204922 -74
rect 204864 -130 204872 -96
rect 204906 -130 204922 -96
rect 204864 -146 204922 -130
rect 202616 -542 202694 -498
rect 202616 -594 202630 -542
rect 202682 -594 202694 -542
rect 202616 -630 202694 -594
rect 173130 -2778 173208 -2732
rect 179394 -2750 179458 -2688
rect 173130 -2812 173156 -2778
rect 173190 -2812 173208 -2778
rect 166558 -2848 166630 -2818
rect 166558 -2882 166573 -2848
rect 166607 -2882 166630 -2848
rect 166558 -2900 166630 -2882
rect 169622 -2870 169682 -2854
rect 166566 -4328 166594 -2900
rect 169622 -2904 169637 -2870
rect 169671 -2904 169682 -2870
rect 169622 -2918 169682 -2904
rect 169624 -3632 169678 -2918
rect 169616 -3652 169692 -3632
rect 169616 -3686 169633 -3652
rect 169667 -3686 169692 -3652
rect 169616 -3702 169692 -3686
rect 173130 -3690 173208 -2812
rect 173130 -3724 173158 -3690
rect 173192 -3724 173208 -3690
rect 173130 -3798 173208 -3724
rect 176548 -2780 176624 -2754
rect 176548 -2814 176569 -2780
rect 176603 -2814 176624 -2780
rect 176548 -3690 176624 -2814
rect 176548 -3724 176567 -3690
rect 176601 -3724 176624 -3690
rect 176548 -3750 176624 -3724
rect 179394 -2784 179412 -2750
rect 179446 -2784 179458 -2750
rect 179394 -3712 179458 -2784
rect 182742 -2804 182784 -2796
rect 182740 -2812 182788 -2804
rect 182738 -2816 182788 -2812
rect 182738 -2850 182746 -2816
rect 182780 -2850 182788 -2816
rect 191452 -2815 191532 -2770
rect 182738 -2856 182788 -2850
rect 187970 -2850 188048 -2826
rect 182738 -2864 182786 -2856
rect 182742 -3642 182784 -2864
rect 187970 -2884 187991 -2850
rect 188025 -2884 188048 -2850
rect 187970 -3608 188048 -2884
rect 191452 -2849 191479 -2815
rect 191513 -2849 191532 -2815
rect 191452 -3223 191532 -2849
rect 195660 -2862 195744 -2816
rect 195660 -2896 195690 -2862
rect 195724 -2896 195744 -2862
rect 195660 -3104 195744 -2896
rect 195660 -3138 195686 -3104
rect 195720 -3138 195744 -3104
rect 195660 -3160 195744 -3138
rect 191452 -3257 191467 -3223
rect 191501 -3257 191532 -3223
rect 191452 -3284 191532 -3257
rect 187970 -3642 187991 -3608
rect 188025 -3642 188048 -3608
rect 182742 -3650 182792 -3642
rect 182742 -3684 182748 -3650
rect 182782 -3684 182792 -3650
rect 187970 -3666 188048 -3642
rect 182742 -3694 182792 -3684
rect 182742 -3704 182784 -3694
rect 179394 -3746 179412 -3712
rect 179446 -3746 179458 -3712
rect 179394 -3782 179458 -3746
rect 166566 -4452 166602 -4328
rect 166560 -4454 166606 -4452
rect 166550 -4460 166618 -4454
rect 166550 -4490 166567 -4460
rect 166552 -4494 166567 -4490
rect 166601 -4494 166618 -4460
rect 166552 -4506 166618 -4494
rect 169618 -4752 169678 -4736
rect 169618 -4786 169635 -4752
rect 169669 -4786 169678 -4752
rect 169618 -4794 169678 -4786
rect 169624 -4942 169676 -4794
rect 169624 -4944 169684 -4942
rect 169622 -4955 169684 -4944
rect 169622 -4989 169636 -4955
rect 169670 -4989 169684 -4955
rect 169622 -5006 169684 -4989
rect 173128 -5604 173204 -5190
rect 176546 -6294 176622 -6246
rect 176546 -6328 176563 -6294
rect 176597 -6328 176622 -6294
rect 176546 -6730 176622 -6328
rect 176546 -6763 176626 -6730
rect 176546 -6797 176572 -6763
rect 176606 -6797 176626 -6763
rect 176546 -6816 176626 -6797
rect 176548 -6820 176626 -6816
rect 179400 -9612 179468 -9590
rect 179400 -9646 179418 -9612
rect 179452 -9646 179468 -9612
rect 179400 -9830 179468 -9646
rect 179400 -9844 179470 -9830
rect 179400 -9878 179420 -9844
rect 179454 -9878 179470 -9844
rect 179400 -9896 179470 -9878
rect 182750 -14818 182810 -14804
rect 182748 -14852 182762 -14818
rect 182796 -14852 182810 -14818
rect 182748 -14862 182810 -14852
rect 182748 -15050 182800 -14862
rect 182742 -15062 182802 -15050
rect 182742 -15096 182752 -15062
rect 182786 -15096 182802 -15062
rect 182742 -15108 182802 -15096
<< via1 >>
rect 203361 178 203413 230
rect 202630 -594 202682 -542
<< metal2 >>
rect 196108 28170 196194 28938
rect 196108 27644 196198 28170
rect 167888 -2118 168006 -2108
rect 196120 -2118 196198 27644
rect 203350 322 203432 332
rect 203348 315 203432 322
rect 203348 259 203363 315
rect 203419 259 203432 315
rect 203348 242 203432 259
rect 203348 230 203420 242
rect 203348 178 203361 230
rect 203413 178 203420 230
rect 203348 164 203420 178
rect 202496 -530 202556 -522
rect 202496 -542 202688 -530
rect 202496 -594 202630 -542
rect 202682 -594 202688 -542
rect 202496 -600 202688 -594
rect 202496 -2118 202556 -600
rect 167888 -2198 202556 -2118
rect 167888 -3814 168006 -2198
rect 196120 -2220 196198 -2198
<< via2 >>
rect 203363 259 203419 315
<< metal3 >>
rect 203346 435 203422 468
rect 203346 378 203354 435
rect 203348 371 203354 378
rect 203418 424 203422 435
rect 203418 371 203430 424
rect 203348 336 203430 371
rect 203350 315 203430 336
rect 203350 259 203363 315
rect 203419 259 203430 315
rect 203350 242 203430 259
<< via3 >>
rect 203354 371 203418 435
<< metal4 >>
rect 201162 31044 201518 31050
rect 197054 30978 201640 31044
rect 201162 30968 201640 30978
rect 201540 25428 201640 30968
rect 201540 25220 201734 25428
rect 201542 648 201734 25220
rect 201542 576 203420 648
rect 201554 414 201720 576
rect 203348 516 203420 576
rect 203346 496 203420 516
rect 203346 435 203422 496
rect 201554 314 201724 414
rect 203346 371 203354 435
rect 203418 424 203422 435
rect 203418 371 203434 424
rect 203346 352 203434 371
rect 166934 -1628 167402 -1624
rect 201558 -1628 201724 314
rect 166934 -1828 201724 -1628
rect 166946 -2842 167064 -1828
rect 166936 -2912 167064 -2842
rect 166936 -4012 167054 -2912
use 9bitdac_layout  9bitdac_layout_0
timestamp 1624221218
transform 1 0 0 0 1 1976
box 0 -1976 198772 52794
use 9bitdac_layout  9bitdac_layout_1
timestamp 1624221218
transform 1 0 -428 0 1 -55716
box 0 -1976 198772 52794
use switch_layout  switch_layout_0
timestamp 1624221218
transform 1 0 202454 0 1 -818
box 40 172 2460 1180
use res250_layout  res250_layout_0
timestamp 1624221218
transform 1 0 165760 0 1 5268
box 218 -342 484 -90
<< labels >>
rlabel locali s 166002 5196 166002 5196 4 x1_vref5
rlabel locali s 166178 4858 166178 4858 4 x2_vref1
rlabel locali s 165594 -52506 165594 -52506 4 inp2
rlabel locali s 830 53968 830 53968 4 inp1
rlabel locali s 202424 -280 202424 -280 4 d9
rlabel locali s 204962 -118 204962 -118 4 out_v
rlabel metal2 s 202538 -566 202538 -566 4 gnd!
rlabel metal4 s 203376 488 203376 488 4 vdd!
rlabel locali s 204708 432 204708 432 4 x1_out_v
rlabel locali s 204730 -712 204730 -712 4 x2_out_v
rlabel locali s 166580 414 166580 414 4 d0
rlabel locali s 169642 144 169642 144 4 d1
rlabel locali s 173170 -566 173170 -566 4 d2
rlabel locali s 176582 -860 176582 -860 4 d3
rlabel locali s 179432 -344 179432 -344 4 d4
rlabel locali s 182764 -170 182764 -170 4 d5
rlabel locali s 188000 -138 188000 -138 4 d6
rlabel locali s 191500 -950 191500 -950 4 d7
rlabel locali s 195706 -1220 195706 -1220 4 d8
<< end >>
