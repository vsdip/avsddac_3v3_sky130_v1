magic
tech sky130A
magscale 1 2
timestamp 1625518311
<< locali >>
rect 236 11484 292 11620
rect 13494 6278 16080 6312
rect 13494 6276 16078 6278
rect 10824 6080 11014 6204
rect 10824 4040 10940 6080
rect 10824 4006 10852 4040
rect 10886 4006 10940 4040
rect 10824 3958 10940 4006
rect 7380 2087 7492 3404
rect 7380 2053 7398 2087
rect 7432 2053 7492 2087
rect 7380 2030 7492 2053
rect 10792 2876 10924 2974
rect 10792 2842 10860 2876
rect 10894 2842 10924 2876
rect 10792 2020 10924 2842
rect 16042 2424 16078 6276
rect 16038 2214 16080 2424
rect 16038 2198 16082 2214
rect 3794 1520 3936 1620
rect 3794 1080 3884 1520
rect 3794 1046 3809 1080
rect 3843 1046 3884 1080
rect 3794 1020 3884 1046
rect 7312 1373 7464 1454
rect 7312 1339 7406 1373
rect 7440 1339 7464 1373
rect 806 856 822 866
rect 800 842 822 856
rect 804 828 822 842
rect 754 503 822 828
rect 754 469 778 503
rect 812 469 822 503
rect 754 438 822 469
rect 3794 582 3884 628
rect 3794 548 3817 582
rect 3851 548 3884 582
rect 3794 460 3884 548
rect 766 163 834 178
rect 766 129 776 163
rect 810 129 834 163
rect 14 -164 76 0
rect 766 -187 834 129
rect 3794 44 3892 460
rect 766 -221 786 -187
rect 820 -221 834 -187
rect 766 -250 834 -221
rect 168 -468 228 -402
rect 762 -525 834 -482
rect 762 -559 782 -525
rect 816 -559 834 -525
rect 762 -1038 834 -559
rect 3802 -508 3892 44
rect 7312 -294 7464 1339
rect 3802 -542 3823 -508
rect 3857 -542 3892 -508
rect 3802 -582 3892 -542
rect 3812 -998 3902 -958
rect 3812 -1032 3835 -998
rect 3869 -1032 3902 -998
rect 3812 -1542 3902 -1032
rect 7320 -965 7420 -294
rect 7320 -999 7348 -965
rect 7382 -999 7420 -965
rect 10792 -974 10958 2020
rect 16040 1784 16082 2198
rect 16038 1776 16082 1784
rect 16038 1344 16080 1776
rect 16208 1061 16372 1072
rect 16208 1027 16216 1061
rect 16250 1027 16372 1061
rect 16208 1016 16372 1027
rect 13784 856 13886 946
rect 7320 -1052 7420 -999
rect 7332 -1769 7432 -1706
rect 7332 -1803 7364 -1769
rect 7398 -1803 7432 -1769
rect 7332 -2636 7432 -1803
rect 10826 -1780 10958 -974
rect 16062 -1396 16098 598
rect 10826 -1814 10886 -1780
rect 10920 -1814 10958 -1780
rect 10826 -1928 10958 -1814
rect 10840 -2820 10972 -2706
rect 10840 -2854 10886 -2820
rect 10920 -2854 10972 -2820
rect 10840 -5868 10972 -2854
rect 16044 -3300 16098 -1396
rect 16044 -5290 16080 -3300
rect 16042 -5652 16082 -5290
rect 13412 -5710 16082 -5652
rect 13412 -5714 16074 -5710
rect -54 -12070 4 -11964
<< viali >>
rect 10852 4006 10886 4040
rect 7398 2053 7432 2087
rect 10860 2842 10894 2876
rect 3809 1046 3843 1080
rect 7406 1339 7440 1373
rect 778 469 812 503
rect 3817 548 3851 582
rect 776 129 810 163
rect 786 -221 820 -187
rect 782 -559 816 -525
rect 3823 -542 3857 -508
rect 3835 -1032 3869 -998
rect 7348 -999 7382 -965
rect 16216 1027 16250 1061
rect 7364 -1803 7398 -1769
rect 10886 -1814 10920 -1780
rect 10886 -2854 10920 -2820
<< metal1 >>
rect 10808 4040 10916 4124
rect 10808 4006 10852 4040
rect 10886 4006 10916 4040
rect 10808 2876 10916 4006
rect 10808 2842 10860 2876
rect 10894 2842 10916 2876
rect 10808 2770 10916 2842
rect 7376 2087 7476 2232
rect 7376 2053 7398 2087
rect 7432 2053 7476 2087
rect 7376 1373 7476 2053
rect 7376 1339 7406 1373
rect 7440 1339 7476 1373
rect 7376 1302 7476 1339
rect 14674 1390 14798 1416
rect 14674 1338 14725 1390
rect 14777 1338 14798 1390
rect 14674 1320 14798 1338
rect 3794 1080 3884 1102
rect 3794 1046 3809 1080
rect 3843 1046 3884 1080
rect 3794 582 3884 1046
rect 16214 1061 16252 1064
rect 16214 1027 16216 1061
rect 16250 1027 16252 1061
rect 16214 1024 16252 1027
rect 16258 1020 16270 1066
rect 16214 1018 16258 1020
rect 3794 548 3817 582
rect 3851 548 3884 582
rect 762 503 830 534
rect 3794 518 3884 548
rect 13936 598 14048 664
rect 13936 546 13952 598
rect 14004 546 14048 598
rect 13936 520 14048 546
rect 762 469 778 503
rect 812 469 830 503
rect 762 163 830 469
rect 762 129 776 163
rect 810 129 830 163
rect 762 106 830 129
rect 762 -187 830 -172
rect 762 -221 786 -187
rect 820 -221 830 -187
rect 762 -525 830 -221
rect 762 -559 782 -525
rect 816 -559 830 -525
rect 762 -600 830 -559
rect 3802 -508 3892 -482
rect 3802 -542 3823 -508
rect 3857 -542 3892 -508
rect 3802 -998 3892 -542
rect 3802 -1032 3835 -998
rect 3869 -1032 3892 -998
rect 3802 -1066 3892 -1032
rect 7328 -965 7428 -912
rect 7328 -999 7348 -965
rect 7382 -999 7428 -965
rect 7328 -1769 7428 -999
rect 7328 -1803 7364 -1769
rect 7398 -1803 7428 -1769
rect 7328 -1842 7428 -1803
rect 10848 -1780 10956 -1624
rect 10848 -1814 10886 -1780
rect 10920 -1814 10956 -1780
rect 10848 -2820 10956 -1814
rect 10848 -2854 10886 -2820
rect 10920 -2854 10956 -2820
rect 10848 -2978 10956 -2854
<< via1 >>
rect 14725 1338 14777 1390
rect 13952 546 14004 598
<< metal2 >>
rect 10460 4878 10550 5848
rect 10460 4866 13424 4878
rect 10460 4774 13484 4866
rect 13394 570 13484 4774
rect 14702 1514 14802 1530
rect 14700 1510 14802 1514
rect 14700 1454 14725 1510
rect 14781 1454 14802 1510
rect 14700 1418 14802 1454
rect 14700 1390 14800 1418
rect 14700 1338 14725 1390
rect 14777 1338 14800 1390
rect 14700 1322 14800 1338
rect 13938 598 14010 632
rect 13938 570 13952 598
rect 13390 546 13952 570
rect 14004 546 14010 598
rect 13390 518 14010 546
rect 13394 -172 13484 518
rect 13388 -254 13484 -172
rect 13388 -4702 13478 -254
rect 13388 -4746 13484 -4702
rect 10758 -6932 10840 -6150
rect 10744 -6936 12360 -6932
rect 13394 -6936 13484 -4746
rect 10744 -7006 13486 -6936
rect 10758 -7010 10840 -7006
rect 12108 -7010 13486 -7006
rect 13394 -7022 13484 -7010
<< via2 >>
rect 14725 1454 14781 1510
<< metal3 >>
rect 14698 1626 14816 1660
rect 14698 1562 14728 1626
rect 14792 1562 14816 1626
rect 14698 1540 14816 1562
rect 14702 1510 14798 1540
rect 14702 1454 14725 1510
rect 14781 1454 14798 1510
rect 14702 1434 14798 1454
<< via3 >>
rect 14728 1562 14792 1626
<< metal4 >>
rect 10134 3322 10222 7012
rect 10134 1824 10224 3322
rect 14698 1824 14814 1828
rect 10130 1712 14814 1824
rect 10134 -5100 10224 1712
rect 14698 1626 14814 1712
rect 14698 1562 14728 1626
rect 14792 1562 14814 1626
rect 14698 1540 14814 1562
use 4bitdac_layout  4bitdac_layout_0
timestamp 1625518311
transform 1 0 -64 0 1 -5936
box -6 -6048 13514 5724
use 4bitdac_layout  4bitdac_layout_1
timestamp 1625518311
transform 1 0 6 0 1 6048
box -6 -6048 13514 5724
use res250_layout  res250_layout_0
timestamp 1625518311
transform 1 0 -230 0 1 -62
box 218 -342 484 -90
use switch_layout  switch_layout_0
timestamp 1625518311
transform 1 0 13800 0 1 336
box 40 154 2460 1180
<< labels >>
rlabel locali s 36 -122 36 -122 4 x1_vref5
rlabel locali s 188 -432 188 -432 4 x2_vref1
rlabel locali s 784 -46 784 -46 4 d0
rlabel locali s 3842 -18 3842 -18 4 d1
rlabel locali s 7356 -74 7356 -74 4 d2
rlabel locali s 10878 -158 10878 -158 4 d3
rlabel locali s 13812 896 13812 896 4 d4
rlabel locali s 16320 1034 16320 1034 4 out_v
rlabel locali s 13596 -5688 13596 -5688 4 x2_out_v
rlabel locali s 13732 6288 13732 6288 4 x1_out_v
rlabel locali s 262 11508 262 11508 4 inp1
rlabel locali s 258 11576 258 11576 4 inp1
rlabel locali s -36 -12014 -36 -12014 4 inp2
rlabel metal4 s 14500 1778 14500 1778 4 vdd!
rlabel metal2 s 13440 532 13440 532 4 gnd!
<< end >>
