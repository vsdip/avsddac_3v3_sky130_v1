magic
tech sky130A
magscale 1 2
timestamp 1640022418
<< locali >>
rect 19916 48682 19962 48686
rect 19916 48680 19964 48682
rect 19916 48672 19966 48680
rect 19916 48638 19924 48672
rect 19958 48670 19966 48672
rect 43760 48670 45162 48678
rect 19958 48640 45162 48670
rect 19958 48638 43838 48640
rect 19916 48632 43838 48638
rect 19916 48630 27254 48632
rect 45116 48624 45162 48640
rect 11768 48096 20162 48100
rect -252 48050 20860 48096
rect -252 48046 11818 48050
rect -252 48040 3448 48046
rect -246 -164 -194 48040
rect 544 47846 602 48006
rect 19916 47982 19976 47990
rect 19916 47948 19930 47982
rect 19964 47948 19976 47982
rect 19916 47940 19976 47948
rect 19918 30780 19964 47940
rect 20810 47820 20858 48050
rect 45116 46140 45166 48624
rect 19918 30744 19970 30780
rect 19922 27384 19970 30744
rect 19916 27342 19970 27384
rect 19916 26696 19964 27342
rect 19916 26662 19966 26696
rect 19918 26004 19966 26662
rect 45116 26240 45170 46140
rect 45116 26204 45180 26240
rect 19918 25974 19970 26004
rect 19922 24586 19970 25974
rect 45120 25704 45180 26204
rect 45122 25350 45176 25704
rect 45316 25065 45562 25086
rect 45316 25031 45340 25065
rect 45374 25031 45562 25065
rect 45316 25018 45562 25031
rect 42884 24848 42968 24952
rect 41604 24610 42370 24614
rect 40178 24554 42372 24610
rect 40178 24550 41694 24554
rect 17260 13452 17380 24516
rect 17260 13418 17300 13452
rect 17334 13418 17380 13452
rect 17260 13380 17380 13418
rect 37596 13344 37638 24484
rect 42332 24162 42372 24554
rect 45176 24166 45216 24602
rect 43884 24162 45222 24166
rect 42332 24122 45222 24162
rect 42332 24120 44692 24122
rect 42332 24116 43924 24120
rect 37596 13310 37602 13344
rect 37636 13310 37638 13344
rect 37596 13294 37638 13310
rect 13936 12996 14044 13104
rect 17230 13014 17360 13046
rect 13946 9290 14034 12996
rect 17230 12980 17280 13014
rect 17314 12980 17360 13014
rect 17230 11702 17360 12980
rect 17230 11514 17368 11702
rect 13928 8130 14034 9290
rect 13928 7460 14016 8130
rect 13928 6810 14024 7460
rect 13928 6776 13962 6810
rect 13996 6776 14024 6810
rect 13930 6740 14024 6776
rect 10834 6284 11118 6382
rect 10838 5450 10908 6284
rect 10830 5384 10908 5450
rect 13928 6216 14016 6278
rect 13928 6182 13952 6216
rect 13986 6182 14016 6216
rect 10830 4776 10904 5384
rect 10824 4474 10904 4776
rect 10824 3867 10898 4474
rect 13928 4124 14016 6182
rect 13930 4052 14012 4124
rect 13930 3918 14042 4052
rect 10824 3833 10845 3867
rect 10879 3833 10898 3867
rect 10824 3800 10898 3833
rect 7484 3468 7582 3552
rect 10812 3531 10886 3560
rect 10812 3497 10819 3531
rect 10853 3497 10886 3531
rect 7486 2912 7540 3468
rect 7482 2115 7542 2912
rect 10812 2874 10886 3497
rect 7482 2081 7493 2115
rect 7527 2081 7542 2115
rect 7482 2030 7542 2081
rect 7482 1739 7542 1760
rect 3982 1706 4008 1724
rect 3982 1202 4040 1706
rect 3982 1168 3995 1202
rect 4029 1168 4040 1202
rect 3982 1154 4040 1168
rect 7482 1705 7493 1739
rect 7527 1705 7542 1739
rect 7482 1074 7542 1705
rect 3970 1012 4044 1022
rect 942 954 1030 980
rect 3970 978 3991 1012
rect 4025 978 4044 1012
rect 942 700 1012 954
rect 3970 930 4044 978
rect 7468 1000 7542 1074
rect 3970 796 4040 930
rect 942 692 1010 700
rect 944 634 1010 692
rect 3966 690 4040 796
rect 944 604 1008 634
rect 936 596 1008 604
rect 3966 600 4020 690
rect 936 562 953 596
rect 987 562 1008 596
rect 936 550 1008 562
rect 944 412 1012 418
rect 944 406 1018 412
rect 944 372 963 406
rect 997 372 1018 406
rect 944 364 1018 372
rect 944 358 1010 364
rect 948 290 1010 358
rect 948 168 1012 290
rect 42 -2 214 34
rect 42 -118 104 -2
rect 944 -28 1012 168
rect 3938 76 4020 600
rect 7468 392 7538 1000
rect 10810 394 10898 2874
rect 13934 1138 14042 3918
rect 17248 1390 17368 11514
rect 34244 7424 34288 13136
rect 37590 12930 37634 12962
rect 37590 12896 37596 12930
rect 37630 12896 37634 12930
rect 37590 12880 37634 12896
rect 34236 7310 34288 7424
rect 34236 6627 34286 7310
rect 34236 6593 34242 6627
rect 34276 6593 34286 6627
rect 34236 6578 34286 6593
rect 31008 6268 31386 6392
rect 31008 6160 31132 6268
rect 34242 6230 34286 6238
rect 34238 6224 34286 6230
rect 34238 6190 34242 6224
rect 34276 6190 34286 6224
rect 34238 6172 34286 6190
rect 31018 4026 31130 6160
rect 31002 3834 31144 4026
rect 31002 3800 31064 3834
rect 31098 3800 31144 3834
rect 31002 3734 31144 3800
rect 27776 2084 27854 3514
rect 27776 2050 27803 2084
rect 27837 2050 27854 2084
rect 27776 1984 27854 2050
rect 31040 3402 31128 3448
rect 31040 3368 31070 3402
rect 31104 3368 31128 3402
rect 3938 38 4018 76
rect -246 -360 -192 -164
rect -246 -362 172 -360
rect 214 -362 308 -350
rect -246 -416 308 -362
rect -118 -418 308 -416
rect 214 -420 308 -418
rect 936 -1568 1012 -28
rect 936 -1940 1014 -1568
rect 936 -2396 1016 -1940
rect 3930 -2024 4018 38
rect 7436 -1950 7548 392
rect 10804 -1788 10898 394
rect 13890 764 14042 1138
rect 13890 -1484 14012 764
rect 17228 -1042 17408 1390
rect 24250 1239 24336 1754
rect 24250 1205 24282 1239
rect 24316 1205 24336 1239
rect 24250 1178 24336 1205
rect 27766 1612 27844 1676
rect 27766 1578 27785 1612
rect 27819 1578 27844 1612
rect 21198 568 21264 920
rect 21198 534 21207 568
rect 21241 534 21264 568
rect 21198 528 21264 534
rect 24238 915 24324 984
rect 24238 881 24270 915
rect 24304 881 24324 915
rect 21206 526 21242 528
rect 21190 358 21256 374
rect 21190 324 21207 358
rect 21241 324 21256 358
rect 21190 68 21256 324
rect 21190 -18 21258 68
rect 20414 -128 20468 -28
rect 21212 -952 21258 -18
rect 24238 -60 24324 881
rect 27766 272 27844 1578
rect 31040 1532 31128 3368
rect 31032 966 31146 1532
rect 31032 516 31176 966
rect 27712 146 27844 272
rect 24238 -912 24298 -60
rect 24236 -929 24298 -912
rect 21206 -966 21268 -952
rect 21206 -1000 21216 -966
rect 21250 -1000 21268 -966
rect 24236 -963 24252 -929
rect 24286 -963 24298 -929
rect 27712 -892 27810 146
rect 27712 -926 27733 -892
rect 27767 -926 27810 -892
rect 27712 -962 27810 -926
rect 31048 -855 31176 516
rect 34242 472 34286 6172
rect 37592 2112 37634 12880
rect 34202 418 34286 472
rect 34202 334 34296 418
rect 34210 -218 34296 334
rect 31048 -889 31101 -855
rect 31135 -889 31176 -855
rect 24236 -996 24298 -963
rect 31048 -978 31176 -889
rect 34202 -318 34296 -218
rect 34202 -902 34288 -318
rect 34202 -936 34220 -902
rect 34254 -936 34288 -902
rect 34202 -954 34288 -936
rect 21206 -1006 21268 -1000
rect 37532 -1042 37652 2112
rect 17198 -1200 37654 -1042
rect 17198 -1216 19098 -1200
rect 27596 -1222 37654 -1200
rect 27596 -1252 31946 -1222
rect 33618 -1470 34274 -1452
rect 20416 -1484 34274 -1470
rect 13890 -1486 34274 -1484
rect 13890 -1520 34224 -1486
rect 34258 -1520 34274 -1486
rect 13890 -1606 34274 -1520
rect 13890 -1620 20582 -1606
rect 33618 -1620 34274 -1606
rect 28184 -1740 31172 -1726
rect 21244 -1756 31172 -1740
rect 14370 -1767 31172 -1756
rect 14370 -1788 31081 -1767
rect 10804 -1801 31081 -1788
rect 31115 -1801 31172 -1767
rect 10804 -1854 31172 -1801
rect 10804 -1868 28408 -1854
rect 10804 -1884 21406 -1868
rect 10804 -1908 14418 -1884
rect 10892 -1916 14418 -1908
rect 7412 -1986 7552 -1950
rect 11356 -1984 11698 -1976
rect 11356 -1986 24578 -1984
rect 7412 -2020 24578 -1986
rect 3930 -2272 4010 -2024
rect 7412 -2052 27818 -2020
rect 7412 -2086 27749 -2052
rect 27783 -2086 27818 -2052
rect 7412 -2120 27818 -2086
rect 7412 -2124 24578 -2120
rect 7412 -2130 11500 -2124
rect 7412 -2148 7552 -2130
rect 3928 -2276 4048 -2272
rect 12266 -2276 20764 -2260
rect 3928 -2285 24300 -2276
rect 3928 -2319 24254 -2285
rect 24288 -2319 24300 -2285
rect 3928 -2342 24300 -2319
rect 3928 -2358 12398 -2342
rect 942 -2398 1016 -2396
rect 21200 -2398 21260 -2390
rect 942 -2400 4086 -2398
rect 19604 -2400 21260 -2398
rect 942 -2405 21260 -2400
rect 942 -2439 21211 -2405
rect 21245 -2439 21260 -2405
rect 942 -2448 21260 -2439
rect 942 -2454 19742 -2448
rect 21200 -2452 21260 -2448
rect 942 -2456 1016 -2454
rect 4060 -2456 19742 -2454
<< viali >>
rect 19924 48638 19958 48672
rect 19930 47948 19964 47982
rect 45340 25031 45374 25065
rect 17300 13418 17334 13452
rect 37602 13310 37636 13344
rect 17280 12980 17314 13014
rect 13962 6776 13996 6810
rect 13952 6182 13986 6216
rect 10845 3833 10879 3867
rect 10819 3497 10853 3531
rect 7493 2081 7527 2115
rect 3995 1168 4029 1202
rect 7493 1705 7527 1739
rect 3991 978 4025 1012
rect 953 562 987 596
rect 963 372 997 406
rect 37596 12896 37630 12930
rect 34242 6593 34276 6627
rect 34242 6190 34276 6224
rect 31064 3800 31098 3834
rect 27803 2050 27837 2084
rect 31070 3368 31104 3402
rect 24282 1205 24316 1239
rect 27785 1578 27819 1612
rect 21207 534 21241 568
rect 24270 881 24304 915
rect 21207 324 21241 358
rect 21216 -1000 21250 -966
rect 24252 -963 24286 -929
rect 27733 -926 27767 -892
rect 31101 -889 31135 -855
rect 34220 -936 34254 -902
rect 34224 -1520 34258 -1486
rect 31081 -1801 31115 -1767
rect 27749 -2086 27783 -2052
rect 24254 -2319 24288 -2285
rect 21211 -2439 21245 -2405
<< metal1 >>
rect 19916 48680 19962 48686
rect 19916 48672 19966 48680
rect 19916 48638 19924 48672
rect 19958 48638 19966 48672
rect 19916 48630 19966 48638
rect 19916 47990 19962 48630
rect 19916 47982 19976 47990
rect 19916 47948 19930 47982
rect 19964 47948 19976 47982
rect 19916 47940 19976 47948
rect 43774 25378 43882 25392
rect 43774 25326 43811 25378
rect 43863 25326 43882 25378
rect 43774 25316 43882 25326
rect 45316 25065 45392 25084
rect 45316 25031 45340 25065
rect 45374 25031 45392 25065
rect 45316 25018 45392 25031
rect 43050 24608 43134 24662
rect 43050 24556 43063 24608
rect 43115 24556 43134 24608
rect 43050 24518 43134 24556
rect 17230 13452 17378 13492
rect 17230 13418 17300 13452
rect 17334 13418 17378 13452
rect 17230 13014 17378 13418
rect 17230 12980 17280 13014
rect 17314 12980 17378 13014
rect 17230 12934 17378 12980
rect 37590 13344 37642 13364
rect 37590 13310 37602 13344
rect 37636 13310 37642 13344
rect 37590 12930 37642 13310
rect 37590 12896 37596 12930
rect 37630 12896 37642 12930
rect 37590 12878 37642 12896
rect 13926 6810 14020 6856
rect 13926 6776 13962 6810
rect 13996 6776 14020 6810
rect 13926 6216 14020 6776
rect 13926 6182 13952 6216
rect 13986 6182 14020 6216
rect 13926 6136 14020 6182
rect 34236 6627 34284 6668
rect 34236 6593 34242 6627
rect 34276 6593 34284 6627
rect 34236 6224 34284 6593
rect 34236 6190 34242 6224
rect 34276 6190 34284 6224
rect 34236 6170 34284 6190
rect 10802 3867 10888 3910
rect 10802 3833 10845 3867
rect 10879 3833 10888 3867
rect 10802 3531 10888 3833
rect 10802 3497 10819 3531
rect 10853 3497 10888 3531
rect 10802 3480 10888 3497
rect 31014 3834 31138 3886
rect 31014 3800 31064 3834
rect 31098 3800 31138 3834
rect 31014 3402 31138 3800
rect 31014 3368 31070 3402
rect 31104 3368 31138 3402
rect 31014 3328 31138 3368
rect 7482 2115 7550 2156
rect 7482 2081 7493 2115
rect 7527 2081 7550 2115
rect 7482 1739 7550 2081
rect 7482 1705 7493 1739
rect 7527 1705 7550 1739
rect 7482 1680 7550 1705
rect 27766 2084 27854 2172
rect 27766 2050 27803 2084
rect 27837 2050 27854 2084
rect 27766 1612 27854 2050
rect 27766 1578 27785 1612
rect 27819 1578 27854 1612
rect 27766 1544 27854 1578
rect 24220 1239 24328 1312
rect 3970 1202 4040 1226
rect 3970 1168 3995 1202
rect 4029 1168 4040 1202
rect 3970 1012 4040 1168
rect 3970 978 3991 1012
rect 4025 978 4040 1012
rect 3970 964 4040 978
rect 24220 1205 24282 1239
rect 24316 1205 24328 1239
rect 24220 915 24328 1205
rect 24220 881 24270 915
rect 24304 881 24328 915
rect 24220 856 24328 881
rect 944 604 1008 614
rect 936 596 1008 604
rect 936 562 953 596
rect 987 562 1008 596
rect 936 526 1008 562
rect 21188 568 21262 592
rect 21188 534 21207 568
rect 21241 534 21262 568
rect 936 518 1010 526
rect 932 474 1020 518
rect 932 470 1012 474
rect 950 424 1012 470
rect 944 412 1012 424
rect 944 406 1018 412
rect 944 372 963 406
rect 997 372 1018 406
rect 944 364 1018 372
rect 944 362 1010 364
rect 21188 358 21262 534
rect 21188 324 21207 358
rect 21241 324 21262 358
rect 21188 312 21262 324
rect 21188 306 21260 312
rect 27712 -884 27808 -828
rect 31048 -855 31176 -802
rect 27712 -892 27812 -884
rect 24236 -929 24298 -892
rect 21206 -966 21268 -952
rect 21206 -1000 21216 -966
rect 21250 -1000 21268 -966
rect 21206 -1006 21268 -1000
rect 24236 -963 24252 -929
rect 24286 -963 24298 -929
rect 27712 -926 27733 -892
rect 27767 -926 27812 -892
rect 27712 -962 27812 -926
rect 21208 -2390 21244 -1006
rect 24236 -2285 24298 -963
rect 27714 -2052 27812 -962
rect 31048 -889 31101 -855
rect 31135 -889 31176 -855
rect 31048 -1658 31176 -889
rect 34194 -902 34280 -876
rect 34194 -936 34220 -902
rect 34254 -936 34280 -902
rect 34194 -1486 34280 -936
rect 34194 -1520 34224 -1486
rect 34258 -1520 34280 -1486
rect 34194 -1612 34280 -1520
rect 31048 -1767 31172 -1658
rect 31048 -1801 31081 -1767
rect 31115 -1801 31172 -1767
rect 31048 -1854 31172 -1801
rect 27714 -2086 27749 -2052
rect 27783 -2086 27812 -2052
rect 27714 -2118 27812 -2086
rect 24236 -2319 24254 -2285
rect 24288 -2319 24298 -2285
rect 24236 -2326 24298 -2319
rect 24242 -2346 24298 -2326
rect 21200 -2405 21260 -2390
rect 21200 -2439 21211 -2405
rect 21245 -2439 21260 -2405
rect 21200 -2452 21260 -2439
<< via1 >>
rect 43811 25326 43863 25378
rect 43063 24556 43115 24608
<< metal2 >>
rect 19138 48464 24104 48470
rect 16350 48460 24104 48464
rect 10768 48384 24104 48460
rect 10768 48378 19186 48384
rect 10768 48374 16396 48378
rect 10768 43598 10832 48374
rect 24060 48362 24104 48384
rect 24060 47762 24116 48362
rect 24060 46508 24126 47762
rect 24060 46470 24132 46508
rect 24066 45216 24132 46470
rect 10768 43518 10854 43598
rect 10778 42020 10854 43518
rect 43792 25464 43886 25482
rect 43792 25408 43809 25464
rect 43865 25408 43886 25464
rect 43792 25378 43886 25408
rect 43792 25326 43811 25378
rect 43863 25326 43886 25378
rect 43792 25316 43886 25326
rect 42950 24620 43128 24624
rect 42944 24608 43128 24620
rect 42944 24556 43063 24608
rect 43115 24556 43128 24608
rect 42944 24526 43128 24556
rect 42944 23834 42980 24526
rect 37200 23790 41970 23802
rect 42944 23790 42976 23834
rect 37200 23756 42976 23790
rect 42944 23754 42976 23756
<< via2 >>
rect 43809 25408 43865 25464
<< metal3 >>
rect 43790 25566 43890 25574
rect 43790 25502 43811 25566
rect 43875 25502 43890 25566
rect 43790 25464 43890 25502
rect 43790 25408 43809 25464
rect 43865 25408 43890 25464
rect 43790 25398 43890 25408
<< via3 >>
rect 43811 25502 43875 25566
<< metal4 >>
rect 7746 48242 7842 48246
rect 22460 48242 22590 48246
rect 7746 48160 22590 48242
rect 7746 47486 7842 48160
rect 22460 48158 22590 48160
rect 22514 47824 22590 48158
rect 38540 26238 42638 26240
rect 43788 26238 43884 26240
rect 38540 26170 43884 26238
rect 38540 26164 42638 26170
rect 43788 25626 43884 26170
rect 43788 25612 43890 25626
rect 43790 25566 43890 25612
rect 43790 25502 43811 25566
rect 43875 25502 43890 25566
rect 43790 25494 43890 25502
use 6bitdac_layout  6bitdac_layout_0
timestamp 1640022418
transform 1 0 244 0 1 24130
box -244 -24130 19716 23842
use 6bitdac_layout  6bitdac_layout_1
timestamp 1640022418
transform 1 0 20506 0 1 24092
box -244 -24130 19716 23842
use res250_layout  res250_layout_0
timestamp 1640022418
transform 1 0 -176 0 1 -20
box 218 -342 484 -90
use switch_layout  switch_layout_0
timestamp 1640022418
transform 1 0 42896 0 1 24336
box 40 154 2460 1180
<< labels >>
rlabel locali s 86 -116 86 -116 4 x1_vref5
rlabel locali s 254 -402 254 -402 4 x2_vref1
rlabel locali s 20436 -88 20436 -88 4 inp2
rlabel locali s 574 47944 574 47944 4 inp1
rlabel locali s 42914 24889 42914 24889 4 d6
rlabel locali s 45424 25060 45424 25060 4 out_v
rlabel metal4 s 43842 25592 43842 25592 4 vdd!
rlabel metal2 s 43000 24558 43000 24558 4 gnd!
rlabel locali s 45196 24296 45196 24296 4 x2_out_v
rlabel locali s 45154 25632 45154 25632 4 x1_out_v
rlabel locali s 978 254 978 254 4 d0
rlabel locali s 3992 214 3992 214 4 d1
rlabel locali s 10852 480 10852 480 4 d3
rlabel locali s 14002 926 14002 926 4 d4
rlabel locali s 17326 810 17326 810 4 d5
rlabel locali s 7486 -1174 7486 -1174 4 d2
<< end >>
