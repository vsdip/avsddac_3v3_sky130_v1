magic
tech sky130A
magscale 1 2
timestamp 1625520517
<< locali >>
rect 45770 51554 90780 51562
rect 95360 51554 96184 51558
rect 45770 51520 96184 51554
rect 45770 51370 45824 51520
rect 95364 51516 96184 51520
rect 45770 51336 45777 51370
rect 45811 51336 45824 51370
rect 45770 51326 45824 51336
rect 96148 51466 96184 51516
rect 21190 51278 21746 51280
rect 21190 51274 37460 51278
rect 20370 51272 37460 51274
rect 20370 51255 48154 51272
rect 20370 51230 20399 51255
rect 20372 51221 20399 51230
rect 20433 51234 48154 51255
rect 20433 51230 21390 51234
rect 20433 51221 20452 51230
rect 20372 51210 20452 51221
rect 45768 51190 45818 51196
rect 45768 51156 45777 51190
rect 45811 51156 45818 51190
rect 796 50625 854 50672
rect 796 50591 811 50625
rect 845 50591 854 50625
rect 796 50586 854 50591
rect 808 50451 844 50452
rect 808 50417 809 50451
rect 843 50417 844 50451
rect 808 50416 844 50417
rect 20382 50411 20456 50432
rect 20382 50377 20399 50411
rect 20433 50377 20456 50411
rect 20382 49560 20456 50377
rect 45768 49816 45818 51156
rect 48098 50662 48154 51234
rect 48092 50643 48158 50662
rect 48092 50609 48111 50643
rect 48145 50609 48158 50643
rect 48092 50594 48158 50609
rect 48098 50590 48154 50594
rect 48114 50441 48158 50446
rect 48114 50407 48119 50441
rect 48153 50407 48158 50441
rect 48114 50402 48158 50407
rect 20380 26192 20460 49560
rect 45768 27474 45816 49816
rect 96148 49202 96190 51466
rect 96146 27622 96190 49202
rect 96146 27580 96196 27622
rect 43122 26731 43162 27404
rect 43122 26697 43124 26731
rect 43158 26697 43162 26731
rect 43122 26682 43162 26697
rect 90376 26755 90468 27392
rect 90376 26721 90401 26755
rect 90435 26721 90468 26755
rect 90376 26658 90468 26721
rect 43110 26517 43164 26526
rect 43110 26483 43120 26517
rect 43154 26483 43164 26517
rect 43110 26472 43164 26483
rect 20380 26162 20466 26192
rect 20386 2810 20466 26162
rect 43116 25406 43164 26472
rect 43110 24386 43164 25406
rect 43102 23928 43164 24386
rect 90376 26401 90434 26460
rect 90376 26367 90389 26401
rect 90423 26367 90434 26401
rect 20386 2312 20472 2810
rect 20382 2288 20472 2312
rect 20382 1880 20468 2288
rect 20600 2184 20702 2358
rect 20776 1880 20878 1974
rect 20382 1790 20884 1880
rect 20386 1788 20884 1790
rect 21292 -1170 21352 48
rect 24370 -1026 24430 192
rect 27710 -818 27770 440
rect 31104 -636 31164 734
rect 34346 -442 34406 1020
rect 37808 -300 37868 1456
rect 43102 1292 43154 23928
rect 67968 2260 68026 2354
rect 43092 -108 43158 1292
rect 48502 39 48572 54
rect 78542 50 78638 662
rect 81690 52 81788 1002
rect 85120 432 85182 1398
rect 85120 98 85190 432
rect 85120 72 85202 98
rect 85126 70 85202 72
rect 48502 5 48523 39
rect 48557 5 48572 39
rect 48502 -10 48572 5
rect 78540 23 78640 50
rect 78540 -11 78570 23
rect 78604 -11 78640 23
rect 81688 16 81790 52
rect 81688 8 81722 16
rect 78540 -38 78640 -11
rect 81690 -18 81722 8
rect 81756 8 81790 16
rect 85126 36 85142 70
rect 85176 36 85202 70
rect 85126 8 85202 36
rect 81756 -18 81788 8
rect 85126 -4 85190 8
rect 78542 -44 78638 -38
rect 81690 -48 81788 -18
rect 88292 -102 89642 -98
rect 90376 -102 90434 26367
rect 93032 26096 93112 27534
rect 96150 27322 96196 27580
rect 96320 27036 96520 27052
rect 96320 27002 96331 27036
rect 96365 27002 96520 27036
rect 96320 26988 96520 27002
rect 93930 26830 93980 26922
rect 96172 26364 96214 26570
rect 96172 26120 96218 26364
rect 96172 26100 96212 26120
rect 93540 26096 96212 26100
rect 93032 26030 96212 26096
rect 93032 26026 93562 26030
rect 88292 -108 90434 -102
rect 43090 -168 90434 -108
rect 43090 -172 85110 -168
rect 85226 -172 90434 -168
rect 43090 -186 43236 -172
rect 88292 -184 90434 -172
rect 85120 -264 85182 -238
rect 85120 -298 85134 -264
rect 85168 -272 85182 -264
rect 85168 -298 85194 -272
rect 37800 -304 63320 -300
rect 85120 -304 85194 -298
rect 37800 -362 85194 -304
rect 37800 -366 85178 -362
rect 37800 -372 63320 -366
rect 37808 -380 37868 -372
rect 34350 -468 34406 -442
rect 81688 -460 81790 -420
rect 44280 -462 81790 -460
rect 44280 -464 81724 -462
rect 39300 -468 81724 -464
rect 34350 -496 81724 -468
rect 81758 -464 81790 -462
rect 81758 -496 81788 -464
rect 34350 -520 81788 -496
rect 34350 -524 81758 -520
rect 34350 -528 70790 -524
rect 34350 -532 44304 -528
rect 34350 -534 39342 -532
rect 34448 -536 39342 -534
rect 31098 -644 36684 -636
rect 42164 -644 57422 -640
rect 31098 -648 65052 -644
rect 31098 -660 72694 -648
rect 78542 -660 78638 -652
rect 31098 -675 78638 -660
rect 31098 -696 78574 -675
rect 31104 -704 31164 -696
rect 36646 -704 78574 -696
rect 42164 -709 78574 -704
rect 78608 -709 78638 -675
rect 42164 -712 78638 -709
rect 57366 -716 78638 -712
rect 65008 -720 78638 -716
rect 78534 -730 78638 -720
rect 27698 -822 33728 -818
rect 27698 -835 75364 -822
rect 27698 -869 75311 -835
rect 75345 -866 75364 -835
rect 75345 -869 75362 -866
rect 27698 -876 75362 -869
rect 27710 -886 27770 -876
rect 75290 -884 75362 -876
rect 71794 -1026 71862 -1022
rect 24370 -1028 71862 -1026
rect 24370 -1062 71812 -1028
rect 71846 -1062 71862 -1028
rect 24370 -1068 58626 -1062
rect 24370 -1070 39590 -1068
rect 71794 -1072 71862 -1062
rect 46996 -1170 48574 -1160
rect 21286 -1172 27752 -1170
rect 40626 -1172 48574 -1170
rect 21286 -1177 48574 -1172
rect 21286 -1211 48521 -1177
rect 48555 -1211 48574 -1177
rect 21286 -1224 48574 -1211
rect 21286 -1230 47092 -1224
rect 21424 -1232 26450 -1230
rect 27734 -1232 40650 -1230
<< viali >>
rect 45777 51336 45811 51370
rect 20399 51221 20433 51255
rect 45777 51156 45811 51190
rect 811 50591 845 50625
rect 809 50417 843 50451
rect 20399 50377 20433 50411
rect 48111 50609 48145 50643
rect 48119 50407 48153 50441
rect 43124 26697 43158 26731
rect 90401 26721 90435 26755
rect 43120 26483 43154 26517
rect 90389 26367 90423 26401
rect 48523 5 48557 39
rect 78570 -11 78604 23
rect 81722 -18 81756 16
rect 85142 36 85176 70
rect 96331 27002 96365 27036
rect 85134 -298 85168 -264
rect 81724 -496 81758 -462
rect 78574 -709 78608 -675
rect 75311 -869 75345 -835
rect 71812 -1062 71846 -1028
rect 48521 -1211 48555 -1177
<< metal1 >>
rect 45766 51372 45824 51384
rect 45764 51370 45824 51372
rect 45764 51336 45777 51370
rect 45811 51336 45824 51370
rect 45764 51326 45824 51336
rect 20376 51255 20450 51276
rect 20376 51221 20399 51255
rect 20433 51221 20450 51255
rect 796 50625 854 50656
rect 796 50591 811 50625
rect 845 50591 854 50625
rect 796 50451 854 50591
rect 796 50417 809 50451
rect 843 50417 854 50451
rect 796 50404 854 50417
rect 20376 50411 20450 51221
rect 45768 51192 45822 51326
rect 45766 51190 45822 51192
rect 45766 51156 45777 51190
rect 45811 51156 45822 51190
rect 45766 51140 45822 51156
rect 48092 50658 48158 50662
rect 48092 50643 48168 50658
rect 48092 50609 48111 50643
rect 48145 50609 48168 50643
rect 48092 50594 48168 50609
rect 48100 50456 48168 50594
rect 20376 50377 20399 50411
rect 20433 50377 20450 50411
rect 48098 50441 48168 50456
rect 48098 50407 48119 50441
rect 48153 50412 48168 50441
rect 48153 50407 48164 50412
rect 48098 50388 48164 50407
rect 20376 50358 20450 50377
rect 94792 27354 94880 27366
rect 94792 27302 94825 27354
rect 94877 27302 94880 27354
rect 94792 27290 94880 27302
rect 96320 27036 96386 27052
rect 96320 27002 96331 27036
rect 96365 27002 96386 27036
rect 96320 26986 96386 27002
rect 43116 26742 43162 26758
rect 90362 26755 90468 26792
rect 43116 26731 43164 26742
rect 43116 26697 43124 26731
rect 43158 26697 43164 26731
rect 43116 26686 43164 26697
rect 90362 26721 90401 26755
rect 90435 26721 90468 26755
rect 43116 26526 43162 26686
rect 43110 26517 43162 26526
rect 43110 26483 43120 26517
rect 43154 26483 43162 26517
rect 43110 26472 43162 26483
rect 43116 26470 43162 26472
rect 90362 26401 90468 26721
rect 94048 26578 94160 26630
rect 94048 26526 94073 26578
rect 94125 26526 94160 26578
rect 94048 26492 94160 26526
rect 90362 26367 90389 26401
rect 90423 26367 90468 26401
rect 90362 26340 90468 26367
rect 48502 46 48572 54
rect 48502 39 48574 46
rect 48502 5 48523 39
rect 48557 5 48574 39
rect 48502 -10 48574 5
rect 48512 -1162 48574 -10
rect 71798 -1022 71858 172
rect 75288 -780 75364 436
rect 85122 98 85186 126
rect 85122 70 85202 98
rect 78540 23 78640 50
rect 78540 -11 78570 23
rect 78604 -11 78640 23
rect 81688 42 81790 52
rect 81688 16 81792 42
rect 81688 8 81722 16
rect 78540 -38 78640 -11
rect 81694 -18 81722 8
rect 81756 -18 81792 16
rect 78542 -675 78638 -38
rect 81694 -462 81792 -18
rect 85122 36 85142 70
rect 85176 36 85202 70
rect 85122 8 85202 36
rect 85122 -206 85186 8
rect 85114 -264 85186 -206
rect 85114 -298 85134 -264
rect 85168 -272 85186 -264
rect 85168 -298 85194 -272
rect 85114 -362 85194 -298
rect 85114 -378 85178 -362
rect 81694 -496 81724 -462
rect 81758 -496 81792 -462
rect 81694 -534 81792 -496
rect 78542 -692 78574 -675
rect 78540 -709 78574 -692
rect 78608 -709 78638 -675
rect 78540 -730 78638 -709
rect 75288 -822 75360 -780
rect 75288 -835 75364 -822
rect 75288 -869 75311 -835
rect 75345 -866 75364 -835
rect 75345 -869 75362 -866
rect 75288 -872 75362 -869
rect 75290 -884 75362 -872
rect 71794 -1028 71862 -1022
rect 71794 -1062 71812 -1028
rect 71846 -1062 71862 -1028
rect 71794 -1072 71862 -1062
rect 48506 -1177 48574 -1162
rect 48506 -1211 48521 -1177
rect 48555 -1211 48574 -1177
rect 48506 -1224 48574 -1211
<< via1 >>
rect 94825 27302 94877 27354
rect 94073 26526 94125 26578
<< metal2 >>
rect 24290 50910 25152 50920
rect 24290 50906 58282 50910
rect 24290 50854 58400 50906
rect 24290 50850 58282 50854
rect 25120 50848 58282 50850
rect 94810 27436 94880 27446
rect 94810 27380 94816 27436
rect 94872 27380 94880 27436
rect 94810 27354 94880 27380
rect 94810 27302 94825 27354
rect 94877 27302 94880 27354
rect 94810 27292 94880 27302
rect 93934 26586 94146 26592
rect 93914 26578 94146 26586
rect 93914 26526 94073 26578
rect 94125 26526 94146 26578
rect 93914 26500 94146 26526
rect 93914 26240 93954 26500
rect 91012 26238 93958 26240
rect 90500 26202 93958 26238
rect 90500 26200 92030 26202
rect 90500 26198 91014 26200
<< via2 >>
rect 94816 27380 94872 27436
<< metal3 >>
rect 94810 27530 94890 27538
rect 94810 27466 94820 27530
rect 94884 27466 94890 27530
rect 94810 27456 94890 27466
rect 94810 27436 94880 27456
rect 94810 27380 94816 27436
rect 94872 27380 94880 27436
rect 94810 27372 94880 27380
<< via3 >>
rect 94820 27466 94884 27530
<< metal4 >>
rect 23762 51496 49764 51500
rect 22752 51434 49764 51496
rect 22752 51432 23808 51434
rect 22764 50622 22848 51432
rect 49692 50314 49762 51434
rect 91334 28070 94890 28140
rect 94816 27590 94890 28070
rect 94810 27584 94890 27590
rect 94810 27530 94888 27584
rect 94810 27466 94820 27530
rect 94884 27466 94888 27530
rect 94810 27460 94888 27466
use switch_layout  switch_layout_0
timestamp 1625520517
transform 1 0 93914 0 1 26310
box 40 154 2460 1180
use 7bitdac_layout  7bitdac_layout_1
timestamp 1625520517
transform 1 0 47558 0 1 2444
box -252 -2456 45562 48686
use 7bitdac_layout  7bitdac_layout_0
timestamp 1625520517
transform 1 0 252 0 1 2456
box -252 -2456 45562 48686
use res250_layout  res250_layout_0
timestamp 1625520517
transform 1 0 20392 0 1 2302
box 218 -342 484 -90
<< labels >>
rlabel locali s 20652 2264 20652 2264 4 x1_vref5
rlabel locali s 20812 1868 20812 1868 4 x2_vref1
rlabel locali s 804 50664 804 50664 4 inp1
rlabel locali s 67994 2294 67994 2294 4 inp2
rlabel locali s 93952 26862 93952 26862 4 d7
rlabel locali s 96452 27014 96452 27014 4 out_v
rlabel locali s 96176 27544 96176 27544 4 x1_out_v
rlabel locali s 96200 26388 96200 26388 4 x2_out_v
rlabel metal2 s 93978 26540 93978 26540 4 gnd!
rlabel metal4 s 94864 27554 94864 27554 4 vdd!
rlabel locali s 43126 44 43126 44 4 d6
rlabel locali s 37842 -218 37842 -218 4 d5
rlabel locali s 34364 612 34364 612 4 d4
rlabel locali s 31132 486 31132 486 4 d3
rlabel locali s 27736 152 27736 152 4 d2
rlabel locali s 24396 40 24396 40 4 d1
rlabel locali s 21316 -64 21316 -64 4 d0
<< end >>
