magic
tech sky130A
magscale 1 2
timestamp 1640022418
<< nwell >>
rect 506 622 602 1172
rect 1210 1100 1380 1122
rect 1166 654 1548 1100
rect 1816 172 2200 624
rect 2010 154 2180 172
<< nmos >>
rect 2010 820 2040 940
rect 1350 340 1380 460
<< pmos >>
rect 1350 700 1380 942
rect 2010 330 2040 570
<< ndiff >>
rect 1920 898 2010 940
rect 1920 864 1938 898
rect 1972 864 2010 898
rect 1920 820 2010 864
rect 2040 898 2130 940
rect 2040 864 2078 898
rect 2112 864 2130 898
rect 2040 820 2130 864
rect 1260 417 1350 460
rect 1260 383 1277 417
rect 1311 383 1350 417
rect 1260 340 1350 383
rect 1380 417 1470 460
rect 1380 383 1418 417
rect 1452 383 1470 417
rect 1380 340 1470 383
<< pdiff >>
rect 1270 868 1350 942
rect 1270 834 1283 868
rect 1317 834 1350 868
rect 1270 800 1350 834
rect 1270 766 1283 800
rect 1317 766 1350 800
rect 1270 700 1350 766
rect 1380 871 1462 942
rect 1380 837 1413 871
rect 1447 837 1462 871
rect 1380 803 1462 837
rect 1380 769 1413 803
rect 1447 769 1462 803
rect 1380 700 1462 769
rect 1930 499 2010 570
rect 1930 465 1943 499
rect 1977 465 2010 499
rect 1930 431 2010 465
rect 1930 397 1943 431
rect 1977 397 2010 431
rect 1930 330 2010 397
rect 2040 501 2122 570
rect 2040 467 2073 501
rect 2107 467 2122 501
rect 2040 433 2122 467
rect 2040 399 2073 433
rect 2107 399 2122 433
rect 2040 330 2122 399
<< ndiffc >>
rect 1938 864 1972 898
rect 2078 864 2112 898
rect 1277 383 1311 417
rect 1418 383 1452 417
<< pdiffc >>
rect 1283 834 1317 868
rect 1283 766 1317 800
rect 1413 837 1447 871
rect 1413 769 1447 803
rect 1943 465 1977 499
rect 1943 397 1977 431
rect 2073 467 2107 501
rect 2073 399 2107 433
<< nsubdiff >>
rect 1246 1057 1334 1086
rect 1246 1023 1273 1057
rect 1307 1023 1334 1057
rect 1246 998 1334 1023
rect 2046 248 2136 276
rect 2046 214 2074 248
rect 2108 214 2136 248
rect 2046 190 2136 214
<< nsubdiffcont >>
rect 1273 1023 1307 1057
rect 2074 214 2108 248
<< poly >>
rect 1350 942 1380 970
rect 2010 940 2040 970
rect 2010 790 2040 820
rect 2170 815 2230 840
rect 2170 790 2183 815
rect 2008 781 2183 790
rect 2217 781 2230 815
rect 2008 760 2230 781
rect 920 580 984 582
rect 730 557 984 580
rect 730 542 935 557
rect 920 523 935 542
rect 969 523 984 557
rect 920 504 984 523
rect 1190 576 1248 582
rect 1350 576 1380 700
rect 1190 557 1380 576
rect 2010 570 2040 760
rect 1190 523 1201 557
rect 1235 540 1380 557
rect 1235 523 1248 540
rect 1190 504 1248 523
rect 1350 460 1380 540
rect 1350 310 1380 340
rect 2010 298 2040 330
<< polycont >>
rect 2183 781 2217 815
rect 935 523 969 557
rect 1201 523 1235 557
<< locali >>
rect 492 992 612 1142
rect 1230 1057 2280 1070
rect 1230 1023 1273 1057
rect 1307 1023 2280 1057
rect 1230 1010 2280 1023
rect 1270 868 1320 1010
rect 1270 834 1283 868
rect 1317 834 1320 868
rect 1270 800 1320 834
rect 1270 766 1283 800
rect 1317 766 1320 800
rect 1270 700 1320 766
rect 1410 871 1462 944
rect 1410 837 1413 871
rect 1447 837 1462 871
rect 1410 803 1462 837
rect 1410 769 1413 803
rect 1447 769 1462 803
rect 842 680 844 682
rect 840 670 870 680
rect 810 667 870 670
rect 810 648 813 667
rect 790 633 813 648
rect 847 633 870 667
rect 790 630 870 633
rect 40 518 196 612
rect 790 610 834 630
rect 840 622 870 630
rect 1410 622 1462 769
rect 1920 898 1980 940
rect 1920 864 1938 898
rect 1972 864 1980 898
rect 1920 730 1980 864
rect 2070 898 2130 1010
rect 2070 864 2078 898
rect 2112 864 2130 898
rect 2070 820 2130 864
rect 2170 830 2230 840
rect 2170 815 2350 830
rect 2170 781 2183 815
rect 2217 813 2350 815
rect 2217 781 2304 813
rect 2170 779 2304 781
rect 2338 779 2350 813
rect 2170 760 2350 779
rect 1408 610 1462 622
rect 1718 726 1980 730
rect 1718 692 1932 726
rect 1966 692 1980 726
rect 1718 678 1980 692
rect 1718 610 1780 678
rect 414 542 570 580
rect 920 557 1248 582
rect 920 523 935 557
rect 969 523 1201 557
rect 1235 523 1248 557
rect 1408 552 1780 610
rect 1408 550 1470 552
rect 1718 550 1780 552
rect 920 504 1248 523
rect 1260 417 1320 460
rect 1260 383 1277 417
rect 1311 383 1320 417
rect 502 192 622 312
rect 1260 260 1320 383
rect 1410 417 1470 550
rect 1410 383 1418 417
rect 1452 383 1470 417
rect 1410 340 1470 383
rect 1930 499 1980 678
rect 1930 465 1943 499
rect 1977 465 1980 499
rect 1930 431 1980 465
rect 1930 397 1943 431
rect 1977 397 1980 431
rect 1930 330 1980 397
rect 2070 501 2122 570
rect 2070 467 2073 501
rect 2107 467 2122 501
rect 2070 433 2122 467
rect 2070 399 2073 433
rect 2107 399 2122 433
rect 2070 260 2122 399
rect 1250 248 2300 260
rect 1250 214 2074 248
rect 2108 214 2300 248
rect 1250 200 2300 214
<< viali >>
rect 813 633 847 667
rect 2304 779 2338 813
rect 1932 692 1966 726
<< metal1 >>
rect 502 980 602 1150
rect 1038 1148 2330 1180
rect 1038 1138 2332 1148
rect 1040 920 1080 1138
rect 920 880 1080 920
rect 920 680 960 880
rect 2292 830 2332 1138
rect 2292 813 2350 830
rect 2292 779 2304 813
rect 2338 779 2350 813
rect 2292 770 2350 779
rect 1920 726 2460 740
rect 1920 692 1932 726
rect 1966 692 2460 726
rect 1920 680 2460 692
rect 790 667 960 680
rect 790 633 813 667
rect 847 633 960 667
rect 790 622 960 633
rect 512 182 612 324
use INV  INV_0
timestamp 1640022418
transform 1 0 602 0 1 622
box -88 -440 290 550
use INV  INV_1
timestamp 1640022418
transform 1 0 224 0 1 622
box -88 -440 290 550
<< labels >>
rlabel metal1 s 544 1068 544 1068 4 vdd!
rlabel metal1 s 540 216 540 216 4 gnd!
rlabel locali s 1576 220 1576 220 4 inp2
rlabel locali s 1778 1032 1778 1032 4 inp1
rlabel locali s 100 566 100 566 4 din
rlabel locali s 470 556 470 556 4 dinb
rlabel poly s 2116 776 2116 776 4 dd
rlabel metal1 s 2112 702 2112 702 4 vout
<< end >>
