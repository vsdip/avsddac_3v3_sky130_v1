magic
tech sky130A
magscale 1 2
timestamp 1624221218
<< checkpaint >>
rect -1348 -1700 1550 1810
<< nwell >>
rect 0 334 288 550
rect 0 0 282 334
<< pwell >>
rect 20 -430 278 -312
<< nmos >>
rect 130 -242 160 -120
<< pmos >>
rect 130 60 160 300
<< ndiff >>
rect 42 -163 130 -120
rect 42 -197 57 -163
rect 91 -197 130 -163
rect 42 -242 130 -197
rect 160 -163 248 -120
rect 160 -197 199 -163
rect 233 -197 248 -163
rect 160 -242 248 -197
<< pdiff >>
rect 50 227 130 300
rect 50 193 63 227
rect 97 193 130 227
rect 50 159 130 193
rect 50 125 63 159
rect 97 125 130 159
rect 50 60 130 125
rect 160 232 242 300
rect 160 198 194 232
rect 228 198 242 232
rect 160 164 242 198
rect 160 130 194 164
rect 228 130 242 164
rect 160 60 242 130
<< ndiffc >>
rect 57 -197 91 -163
rect 199 -197 233 -163
<< pdiffc >>
rect 63 193 97 227
rect 63 125 97 159
rect 194 198 228 232
rect 194 130 228 164
<< psubdiff >>
rect 20 -368 278 -312
rect 20 -402 97 -368
rect 131 -402 179 -368
rect 213 -402 278 -368
rect 20 -430 278 -402
<< nsubdiff >>
rect 40 451 250 498
rect 40 447 166 451
rect 40 413 94 447
rect 128 417 166 447
rect 200 417 250 451
rect 128 413 250 417
rect 40 378 250 413
<< psubdiffcont >>
rect 97 -402 131 -368
rect 179 -402 213 -368
<< nsubdiffcont >>
rect 94 413 128 447
rect 166 417 200 451
<< poly >>
rect 130 300 160 330
rect -88 -39 -30 -10
rect -88 -73 -76 -39
rect -42 -40 -30 -39
rect 130 -40 160 60
rect -42 -73 160 -40
rect -88 -80 160 -73
rect -88 -102 -30 -80
rect 130 -120 160 -80
rect 130 -270 160 -242
<< polycont >>
rect -76 -73 -42 -39
<< locali >>
rect 10 451 270 520
rect 10 447 166 451
rect 10 425 94 447
rect 10 391 41 425
rect 75 413 94 425
rect 128 417 166 447
rect 200 425 270 451
rect 200 417 213 425
rect 128 413 213 417
rect 75 391 213 413
rect 247 391 270 425
rect 10 368 270 391
rect 50 302 100 368
rect 50 227 102 302
rect 50 193 63 227
rect 97 193 102 227
rect 50 159 102 193
rect 50 125 63 159
rect 97 125 102 159
rect 50 58 102 125
rect 190 232 242 300
rect 190 198 194 232
rect 228 198 242 232
rect 190 164 242 198
rect 190 130 194 164
rect 228 130 242 164
rect 190 60 242 130
rect -88 -39 -30 -10
rect -88 -73 -76 -39
rect -42 -73 -30 -39
rect -88 -102 -30 -73
rect 190 -120 240 60
rect 40 -163 100 -120
rect 40 -197 57 -163
rect 91 -197 100 -163
rect 40 -310 100 -197
rect 190 -163 248 -120
rect 190 -197 199 -163
rect 233 -197 248 -163
rect 190 -240 248 -197
rect 20 -336 280 -310
rect 20 -370 52 -336
rect 86 -338 280 -336
rect 86 -368 224 -338
rect 86 -370 97 -368
rect 20 -402 97 -370
rect 131 -402 179 -368
rect 213 -372 224 -368
rect 258 -372 280 -338
rect 213 -402 280 -372
rect 20 -430 280 -402
<< viali >>
rect 41 391 75 425
rect 213 391 247 425
rect 52 -370 86 -336
rect 224 -372 258 -338
<< metal1 >>
rect 0 425 282 528
rect 0 420 41 425
rect -2 391 41 420
rect 75 391 213 425
rect 247 420 282 425
rect 247 391 278 420
rect -2 358 278 391
rect 8 -336 290 -298
rect 8 -370 52 -336
rect 86 -338 290 -336
rect 86 -370 224 -338
rect 8 -372 224 -370
rect 258 -372 290 -338
rect 8 -440 290 -372
<< end >>
