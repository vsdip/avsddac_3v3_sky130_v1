* SPICE3 file created from res_nd_500.ext - technology: sky130A

.option scale=10000u

X0 a_119_n123# a_264_n120# SUB sky130_fd_pr__res_generic_nd w=27 l=124
