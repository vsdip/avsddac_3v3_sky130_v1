* SPICE3 file created from 8bitdac_layout.ext - technology: sky130A

.option scale=10000u

X0 switch_layout_0/dd switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1 switch_layout_0/dd switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2 switch_layout_0/dinb d7 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X3 switch_layout_0/dinb d7 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X4 x1_out_v switch_layout_0/dd out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X5 out_v switch_layout_0/dinb x1_out_v switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X6 x2_out_v switch_layout_0/dd out_v switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X7 out_v switch_layout_0/dinb x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X8 7bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X9 7bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X10 7bitdac_layout_0/switch_layout_0/dinb d6 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X11 7bitdac_layout_0/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X12 7bitdac_layout_0/x1_out_v 7bitdac_layout_0/switch_layout_0/dd x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X13 x1_out_v 7bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/x1_out_v 7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X14 7bitdac_layout_0/x2_out_v 7bitdac_layout_0/switch_layout_0/dd x1_out_v 7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X15 x1_out_v 7bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X16 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X17 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X18 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X19 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X20 7bitdac_layout_0/6bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X21 7bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X22 7bitdac_layout_0/6bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X23 7bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X24 7bitdac_layout_0/6bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X25 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X26 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X27 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X28 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X29 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X30 7bitdac_layout_0/6bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X31 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X32 7bitdac_layout_0/6bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X33 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X34 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X35 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X36 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X37 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X38 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X39 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X40 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X41 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X42 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X43 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X44 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X45 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X46 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X47 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X48 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X49 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X50 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X51 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X52 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X53 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X54 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X55 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X56 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X57 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X58 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X59 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X60 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X61 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X62 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X63 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X64 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X65 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X66 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X67 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X68 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X69 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X70 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X71 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X72 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X73 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X74 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X75 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X76 inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X77 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X78 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X79 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X80 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X81 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X82 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X83 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X84 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X85 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X86 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X87 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X88 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X89 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X90 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X91 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X92 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X93 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X94 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X95 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X96 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X97 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X98 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X99 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X100 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X101 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X102 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X103 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X104 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X105 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X106 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X107 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X108 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X109 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X110 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X111 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X112 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X113 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X114 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X115 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X116 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X117 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X118 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X119 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X120 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X121 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X122 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X123 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X124 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X125 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X126 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X127 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X128 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X129 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X130 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X131 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X132 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X133 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X134 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X135 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X136 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X137 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X138 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X139 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X140 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X141 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X142 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X143 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X144 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X145 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X146 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X147 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X148 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X149 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X150 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X151 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X152 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X153 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X154 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X155 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X156 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X157 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X158 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X159 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X160 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X161 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X162 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X163 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X164 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X165 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X166 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X167 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X168 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X169 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X170 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X171 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X172 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X173 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X174 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X175 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X176 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X177 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X178 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X179 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X180 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X181 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X182 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X183 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X184 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X185 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X186 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X187 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X188 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X189 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X190 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X191 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X192 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X193 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X194 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X195 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X196 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X197 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X198 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X199 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X200 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X201 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X202 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X203 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X204 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X205 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X206 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X207 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X208 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X209 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X210 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X211 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X212 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X213 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X214 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X215 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X216 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X217 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X218 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X219 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X220 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X221 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X222 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X223 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X224 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X225 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X226 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X227 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X228 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X229 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X230 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X231 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X232 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X233 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X234 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X235 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X236 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X237 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X238 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X239 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X240 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X241 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X242 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X243 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X244 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X245 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X246 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X247 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X248 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X249 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X250 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X251 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X252 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X253 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X254 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X255 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X256 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X257 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X258 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X259 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X260 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X261 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X262 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X263 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X264 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X265 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X266 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X267 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X268 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X269 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X270 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X271 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X272 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X273 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X274 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X275 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X276 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X277 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X278 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X279 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X280 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X281 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X282 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X283 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X284 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X285 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X286 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X287 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X288 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X289 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X290 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X291 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X292 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X293 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X294 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X295 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X296 7bitdac_layout_0/6bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X297 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X298 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X299 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X300 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X301 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X302 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X303 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X304 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X305 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X306 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X307 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X308 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X309 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X310 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X311 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X312 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X313 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X314 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X315 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X316 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X317 7bitdac_layout_0/6bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X318 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X319 7bitdac_layout_0/6bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X320 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X321 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X322 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X323 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X324 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X325 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X326 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X327 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X328 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X329 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X330 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X331 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X332 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X333 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X334 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X335 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X336 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X337 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X338 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X339 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X340 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X341 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X342 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X343 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X344 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X345 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X346 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X347 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X348 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X349 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X350 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X351 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X352 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X353 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X354 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X355 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X356 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X357 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X358 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X359 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X360 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X361 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X362 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X363 7bitdac_layout_0/6bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X364 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X365 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X366 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X367 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X368 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X369 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X370 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X371 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X372 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X373 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X374 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X375 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X376 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X377 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X378 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X379 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X380 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X381 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X382 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X383 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X384 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X385 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X386 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X387 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X388 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X389 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X390 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X391 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X392 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X393 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X394 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X395 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X396 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X397 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X398 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X399 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X400 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X401 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X402 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X403 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X404 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X405 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X406 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X407 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X408 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X409 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X410 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X411 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X412 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X413 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X414 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X415 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X416 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X417 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X418 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X419 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X420 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X421 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X422 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X423 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X424 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X425 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X426 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X427 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X428 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X429 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X430 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X431 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X432 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X433 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X434 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X435 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X436 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X437 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X438 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X439 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X440 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X441 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X442 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X443 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X444 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X445 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X446 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X447 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X448 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X449 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X450 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X451 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X452 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X453 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X454 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X455 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X456 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X457 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X458 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X459 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X460 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X461 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X462 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X463 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X464 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X465 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X466 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X467 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X468 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X469 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X470 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X471 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X472 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X473 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X474 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X475 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X476 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X477 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X478 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X479 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X480 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X481 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X482 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X483 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X484 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X485 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X486 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X487 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X488 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X489 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X490 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X491 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X492 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X493 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X494 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X495 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X496 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X497 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X498 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X499 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X500 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X501 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X502 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X503 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X504 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X505 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X506 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X507 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X508 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X509 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X510 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X511 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X512 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X513 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X514 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X515 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X516 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X517 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X518 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X519 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X520 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X521 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X522 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X523 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X524 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X525 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X526 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X527 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X528 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X529 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X530 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X531 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X532 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X533 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X534 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X535 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X536 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X537 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X538 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X539 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X540 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X541 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X542 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X543 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X544 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X545 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X546 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X547 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X548 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X549 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X550 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X551 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X552 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X553 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X554 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X555 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X556 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X557 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X558 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X559 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X560 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X561 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X562 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X563 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X564 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X565 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X566 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X567 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X568 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X569 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X570 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X571 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X572 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X573 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X574 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X575 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X576 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X577 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X578 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X579 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X580 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X581 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X582 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X583 7bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X584 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X585 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X586 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X587 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X588 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X589 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X590 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X591 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X592 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X593 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X594 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X595 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X596 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X597 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X598 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X599 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X600 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X601 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X602 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X603 7bitdac_layout_0/6bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X604 7bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X605 7bitdac_layout_0/6bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X606 7bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X607 7bitdac_layout_0/6bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X608 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X609 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X610 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X611 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X612 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X613 7bitdac_layout_0/6bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X614 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X615 7bitdac_layout_0/6bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X616 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X617 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X618 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X619 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X620 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X621 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X622 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X623 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X624 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X625 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X626 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X627 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X628 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X629 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X630 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X631 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X632 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X633 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X634 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X635 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X636 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X637 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X638 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X639 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X640 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X641 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X642 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X643 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X644 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X645 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X646 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X647 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X648 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X649 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X650 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X651 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X652 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X653 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X654 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X655 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X656 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X657 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X658 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X659 7bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X660 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X661 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X662 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X663 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X664 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X665 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X666 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X667 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X668 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X669 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X670 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X671 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X672 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X673 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X674 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X675 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X676 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X677 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X678 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X679 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X680 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X681 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X682 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X683 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X684 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X685 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X686 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X687 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X688 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X689 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X690 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X691 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X692 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X693 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X694 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X695 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X696 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X697 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X698 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X699 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X700 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X701 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X702 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X703 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X704 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X705 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X706 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X707 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X708 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X709 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X710 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X711 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X712 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X713 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X714 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X715 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X716 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X717 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X718 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X719 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X720 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X721 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X722 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X723 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X724 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X725 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X726 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X727 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X728 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X729 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X730 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X731 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X732 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X733 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X734 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X735 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X736 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X737 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X738 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X739 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X740 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X741 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X742 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X743 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X744 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X745 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X746 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X747 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X748 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X749 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X750 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X751 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X752 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X753 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X754 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X755 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X756 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X757 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X758 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X759 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X760 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X761 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X762 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X763 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X764 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X765 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X766 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X767 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X768 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X769 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X770 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X771 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X772 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X773 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X774 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X775 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X776 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X777 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X778 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X779 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X780 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X781 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X782 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X783 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X784 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X785 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X786 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X787 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X788 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X789 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X790 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X791 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X792 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X793 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X794 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X795 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X796 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X797 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X798 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X799 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X800 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X801 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X802 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X803 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X804 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X805 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X806 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X807 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X808 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X809 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X810 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X811 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X812 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X813 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X814 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X815 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X816 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X817 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X818 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X819 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X820 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X821 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X822 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X823 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X824 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X825 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X826 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X827 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X828 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X829 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X830 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X831 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X832 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X833 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X834 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X835 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X836 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X837 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X838 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X839 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X840 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X841 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X842 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X843 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X844 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X845 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X846 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X847 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X848 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X849 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X850 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X851 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X852 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X853 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X854 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X855 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X856 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X857 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X858 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X859 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X860 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X861 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X862 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X863 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X864 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X865 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X866 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X867 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X868 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X869 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X870 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X871 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X872 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X873 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X874 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X875 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X876 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X877 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X878 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X879 7bitdac_layout_0/6bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X880 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X881 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X882 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X883 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X884 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X885 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X886 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X887 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X888 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X889 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X890 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X891 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X892 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X893 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X894 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X895 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X896 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X897 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X898 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X899 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X900 7bitdac_layout_0/6bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X901 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X902 7bitdac_layout_0/6bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X903 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X904 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X905 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X906 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X907 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X908 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X909 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X910 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X911 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X912 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X913 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X914 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X915 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X916 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X917 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X918 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X919 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X920 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X921 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X922 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X923 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X924 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X925 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X926 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X927 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X928 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X929 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X930 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X931 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X932 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X933 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X934 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X935 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X936 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X937 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X938 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X939 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X940 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X941 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X942 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X943 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X944 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X945 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X946 7bitdac_layout_0/6bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X947 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X948 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X949 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X950 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X951 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X952 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X953 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X954 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X955 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X956 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X957 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X958 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X959 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X960 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X961 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X962 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X963 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X964 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X965 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X966 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X967 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X968 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X969 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X970 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X971 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X972 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X973 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X974 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X975 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X976 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X977 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X978 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X979 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X980 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X981 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X982 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X983 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X984 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X985 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X986 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X987 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X988 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X989 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X990 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X991 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X992 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X993 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X994 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X995 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X996 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X997 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X998 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X999 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1000 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1001 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1002 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1003 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1004 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1005 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1006 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1007 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1008 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1009 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1010 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1011 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1012 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1013 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1014 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1015 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1016 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1017 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1018 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1019 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1020 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1021 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1022 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1023 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1024 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1025 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1026 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1027 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1028 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1029 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1030 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1031 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1032 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1033 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1034 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1035 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1036 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1037 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1038 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1039 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1040 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1041 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1042 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1043 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1044 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1045 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1046 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1047 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1048 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1049 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1050 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1051 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1052 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1053 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1054 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1055 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1056 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1057 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1058 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1059 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1060 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1061 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1062 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1063 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1064 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1065 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1066 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1067 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1068 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1069 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1070 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1071 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1072 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1073 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1074 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1075 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1076 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1077 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1078 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1079 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1080 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1081 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1082 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1083 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1084 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1085 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1086 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1087 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1088 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1089 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1090 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1091 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1092 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1093 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1094 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1095 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1096 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1097 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1098 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1099 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1100 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1101 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1102 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1103 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1104 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1105 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1106 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1107 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1108 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1109 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1110 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1111 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1112 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1113 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1114 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1115 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1116 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1117 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1118 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1119 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1120 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1121 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1122 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1123 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1124 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1125 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1126 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1127 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1128 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1129 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1130 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1131 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1132 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1133 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1134 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1135 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1136 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1137 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1138 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1139 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1140 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1141 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1142 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1143 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1144 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1145 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1146 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1147 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1148 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1149 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1150 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1151 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1152 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1153 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1154 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1155 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1156 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1157 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1158 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1159 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1160 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1161 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1162 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1163 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1164 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1165 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1166 x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1167 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1168 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1169 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1170 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1171 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1172 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1173 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1174 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1175 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1176 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1177 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1178 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1179 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1180 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1181 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1182 7bitdac_layout_0/x1_vref5 7bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1183 7bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1184 7bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1185 7bitdac_layout_1/switch_layout_0/dinb d6 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1186 7bitdac_layout_1/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1187 7bitdac_layout_1/x1_out_v 7bitdac_layout_1/switch_layout_0/dd x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1188 x2_out_v 7bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/x1_out_v 7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1189 7bitdac_layout_1/x2_out_v 7bitdac_layout_1/switch_layout_0/dd x2_out_v 7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1190 x2_out_v 7bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1191 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1192 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1193 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1194 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1195 7bitdac_layout_1/6bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1196 7bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1197 7bitdac_layout_1/6bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1198 7bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1199 7bitdac_layout_1/6bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1200 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1201 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1202 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1203 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1204 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1205 7bitdac_layout_1/6bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1206 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1207 7bitdac_layout_1/6bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1208 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1209 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1210 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1211 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1212 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1213 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1214 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1215 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1216 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1217 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1218 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1219 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1220 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1221 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1222 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1223 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1224 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1225 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1226 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1227 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1228 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1229 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1230 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1231 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1232 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1233 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1234 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1235 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1236 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1237 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1238 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1239 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1240 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1241 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1242 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1243 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1244 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1245 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1246 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1247 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1248 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1249 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1250 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1251 x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1252 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1253 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1254 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1255 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1256 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1257 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1258 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1259 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1260 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1261 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1262 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1263 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1264 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1265 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1266 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1267 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1268 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1269 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1270 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1271 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1272 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1273 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1274 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1275 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1276 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1277 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1278 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1279 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1280 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1281 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1282 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1283 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1284 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1285 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1286 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1287 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1288 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1289 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1290 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1291 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1292 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1293 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1294 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1295 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1296 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1297 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1298 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1299 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1300 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1301 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1302 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1303 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1304 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1305 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1306 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1307 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1308 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1309 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1310 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1311 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1312 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1313 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1314 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1315 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1316 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1317 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1318 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1319 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1320 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1321 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1322 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1323 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1324 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1325 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1326 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1327 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1328 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1329 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1330 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1331 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1332 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1333 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1334 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1335 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1336 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1337 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1338 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1339 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1340 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1341 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1342 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1343 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1344 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1345 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1346 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1347 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1348 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1349 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1350 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1351 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1352 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1353 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1354 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1355 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1356 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1357 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1358 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1359 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1360 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1361 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1362 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1363 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1364 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1365 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1366 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1367 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1368 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1369 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1370 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1371 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1372 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1373 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1374 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1375 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1376 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1377 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1378 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1379 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1380 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1381 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1382 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1383 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1384 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1385 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1386 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1387 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1388 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1389 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1390 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1391 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1392 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1393 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1394 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1395 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1396 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1397 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1398 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1399 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1400 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1401 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1402 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1403 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1404 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1405 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1406 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1407 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1408 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1409 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1410 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1411 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1412 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1413 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1414 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1415 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1416 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1417 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1418 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1419 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1420 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1421 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1422 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1423 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1424 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1425 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1426 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1427 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1428 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1429 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1430 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1431 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1432 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1433 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1434 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1435 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1436 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1437 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1438 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1439 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1440 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1441 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1442 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1443 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1444 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1445 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1446 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1447 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1448 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1449 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1450 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1451 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1452 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1453 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1454 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1455 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1456 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1457 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1458 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1459 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1460 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1461 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1462 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1463 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1464 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1465 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1466 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1467 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1468 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1469 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1470 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1471 7bitdac_layout_1/6bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1472 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1473 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1474 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1475 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1476 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1477 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1478 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1479 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1480 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1481 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1482 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1483 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1484 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1485 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1486 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1487 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1488 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1489 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1490 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1491 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1492 7bitdac_layout_1/6bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1493 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1494 7bitdac_layout_1/6bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1495 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1496 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1497 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1498 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1499 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1500 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1501 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1502 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1503 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1504 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1505 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1506 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1507 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1508 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1509 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1510 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1511 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1512 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1513 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1514 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1515 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1516 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1517 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1518 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1519 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1520 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1521 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1522 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1523 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1524 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1525 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1526 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1527 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1528 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1529 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1530 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1531 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1532 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1533 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1534 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1535 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1536 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1537 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1538 7bitdac_layout_1/6bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1539 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1540 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1541 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1542 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1543 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1544 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1545 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1546 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1547 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1548 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1549 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1550 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1551 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1552 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1553 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1554 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1555 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1556 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1557 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1558 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1559 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1560 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1561 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1562 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1563 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1564 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1565 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1566 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1567 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1568 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1569 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1570 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1571 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1572 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1573 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1574 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1575 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1576 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1577 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1578 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1579 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1580 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1581 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1582 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1583 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1584 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1585 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1586 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1587 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1588 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1589 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1590 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1591 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1592 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1593 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1594 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1595 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1596 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1597 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1598 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1599 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1600 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1601 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1602 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1603 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1604 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1605 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1606 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1607 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1608 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1609 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1610 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1611 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1612 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1613 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1614 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1615 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1616 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1617 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1618 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1619 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1620 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1621 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1622 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1623 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1624 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1625 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1626 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1627 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1628 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1629 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1630 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1631 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1632 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1633 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1634 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1635 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1636 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1637 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1638 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1639 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1640 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1641 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1642 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1643 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1644 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1645 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1646 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1647 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1648 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1649 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1650 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1651 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1652 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1653 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1654 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1655 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1656 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1657 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1658 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1659 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1660 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1661 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1662 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1663 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1664 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1665 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1666 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1667 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1668 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1669 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1670 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1671 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1672 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1673 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1674 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1675 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1676 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1677 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1678 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1679 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1680 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1681 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1682 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1683 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1684 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1685 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1686 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1687 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1688 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1689 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1690 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1691 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1692 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1693 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1694 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1695 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1696 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1697 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1698 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1699 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1700 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1701 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1702 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1703 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1704 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1705 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1706 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1707 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1708 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1709 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1710 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1711 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1712 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1713 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1714 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1715 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1716 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1717 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1718 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1719 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1720 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1721 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1722 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1723 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1724 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1725 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1726 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1727 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1728 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1729 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1730 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1731 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1732 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1733 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1734 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1735 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1736 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1737 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1738 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1739 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1740 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1741 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1742 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1743 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1744 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1745 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1746 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1747 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1748 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1749 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1750 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1751 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1752 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1753 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1754 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1755 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1756 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1757 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1758 7bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1759 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1760 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1761 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1762 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1763 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1764 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1765 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1766 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1767 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1768 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1769 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1770 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1771 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1772 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1773 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1774 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1775 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1776 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1777 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1778 7bitdac_layout_1/6bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1779 7bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1780 7bitdac_layout_1/6bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1781 7bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1782 7bitdac_layout_1/6bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1783 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1784 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1785 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1786 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1787 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1788 7bitdac_layout_1/6bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1789 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1790 7bitdac_layout_1/6bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1791 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1792 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1793 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1794 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1795 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1796 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1797 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1798 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1799 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1800 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1801 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1802 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1803 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1804 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1805 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1806 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1807 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1808 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1809 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1810 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1811 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1812 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1813 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1814 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1815 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1816 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1817 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1818 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1819 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1820 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1821 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1822 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1823 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1824 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1825 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1826 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1827 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1828 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1829 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1830 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1831 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1832 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1833 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1834 7bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1835 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1836 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1837 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1838 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1839 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1840 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1841 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1842 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1843 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1844 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1845 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1846 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1847 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1848 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1849 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1850 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1851 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1852 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1853 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1854 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1855 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1856 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1857 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1858 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1859 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1860 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1861 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1862 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1863 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1864 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1865 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1866 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1867 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1868 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1869 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1870 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1871 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1872 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1873 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1874 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1875 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1876 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1877 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1878 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1879 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1880 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1881 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1882 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1883 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1884 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1885 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1886 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1887 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1888 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1889 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1890 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1891 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1892 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1893 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1894 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1895 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1896 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1897 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1898 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1899 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1900 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1901 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1902 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1903 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1904 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1905 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1906 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1907 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1908 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1909 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1910 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1911 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1912 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1913 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1914 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1915 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1916 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1917 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1918 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1919 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1920 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1921 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1922 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1923 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1924 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1925 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1926 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1927 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1928 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1929 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1930 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1931 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1932 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1933 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1934 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1935 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1936 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1937 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1938 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1939 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1940 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1941 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1942 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1943 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1944 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1945 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1946 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1947 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1948 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1949 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1950 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1951 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1952 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1953 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1954 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1955 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1956 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1957 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1958 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1959 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1960 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1961 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1962 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1963 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1964 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1965 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1966 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1967 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1968 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1969 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1970 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1971 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1972 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1973 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X1974 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X1975 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1976 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1977 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1978 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1979 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1980 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1981 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1982 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1983 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1984 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1985 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1986 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1987 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1988 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1989 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1990 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1991 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1992 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1993 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X1994 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X1995 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1996 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X1997 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X1998 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X1999 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2000 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2001 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2002 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2003 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2004 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2005 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2006 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2007 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2008 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2009 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2010 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2011 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2012 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2013 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2014 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2015 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2016 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2017 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2018 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2019 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2020 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2021 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2022 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2023 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2024 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2025 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2026 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2027 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2028 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2029 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2030 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2031 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2032 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2033 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2034 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2035 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2036 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2037 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2038 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2039 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2040 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2041 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2042 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2043 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2044 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2045 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2046 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2047 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2048 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2049 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2050 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2051 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2052 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2053 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2054 7bitdac_layout_1/6bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2055 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2056 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2057 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2058 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2059 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2060 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2061 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2062 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2063 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2064 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2065 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2066 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2067 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2068 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2069 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2070 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2071 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2072 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2073 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2074 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2075 7bitdac_layout_1/6bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2076 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2077 7bitdac_layout_1/6bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2078 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2079 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2080 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2081 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2082 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2083 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2084 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2085 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2086 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2087 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2088 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2089 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2090 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2091 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2092 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2093 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2094 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2095 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2096 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2097 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2098 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2099 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2100 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2101 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2102 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2103 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2104 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2105 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2106 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2107 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2108 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2109 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2110 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2111 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2112 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2113 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2114 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2115 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2116 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2117 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2118 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2119 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2120 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2121 7bitdac_layout_1/6bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2122 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2123 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2124 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2125 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2126 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2127 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2128 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2129 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2130 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2131 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2132 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2133 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2134 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2135 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2136 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2137 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2138 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2139 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2140 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2141 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2142 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2143 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2144 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2145 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2146 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2147 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2148 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2149 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2150 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2151 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2152 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2153 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2154 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2155 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2156 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2157 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2158 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2159 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2160 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2161 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2162 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2163 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2164 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2165 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2166 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2167 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2168 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2169 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2170 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2171 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2172 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2173 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2174 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2175 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2176 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2177 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2178 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2179 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2180 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2181 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2182 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2183 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2184 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2185 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2186 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2187 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2188 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2189 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2190 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2191 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2192 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2193 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2194 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2195 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2196 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2197 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2198 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2199 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2200 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2201 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2202 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2203 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2204 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2205 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2206 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2207 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2208 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2209 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2210 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2211 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2212 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2213 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2214 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2215 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2216 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2217 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2218 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2219 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2220 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2221 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2222 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2223 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2224 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2225 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2226 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2227 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2228 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2229 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2230 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2231 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2232 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2233 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2234 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2235 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2236 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2237 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2238 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2239 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2240 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2241 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2242 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2243 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2244 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2245 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2246 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2247 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2248 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2249 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2250 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2251 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2252 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2253 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2254 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2255 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2256 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2257 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2258 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2259 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2260 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2261 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2262 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2263 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2264 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2265 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2266 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2267 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2268 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2269 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2270 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2271 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2272 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2273 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2274 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2275 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2276 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2277 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2278 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2279 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2280 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2281 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2282 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2283 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2284 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2285 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2286 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2287 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2288 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2289 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2290 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2291 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2292 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2293 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2294 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2295 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2296 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2297 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2298 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2299 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2300 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2301 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2302 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2303 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2304 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2305 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2306 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2307 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2308 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2309 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2310 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2311 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2312 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2313 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2314 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2315 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2316 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2317 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2318 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2319 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2320 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2321 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2322 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2323 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2324 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2325 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2326 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2327 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2328 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2329 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2330 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2331 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2332 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2333 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2334 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2335 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2336 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2337 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2338 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2339 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2340 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2341 inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2342 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb inp2 gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2343 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2344 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2345 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 gnd gnd sky130_fd_pr__nfet_01v8 w=61 l=15
X2346 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=120 l=15
X2347 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2348 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=121 l=15
X2349 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=120 l=15
X2350 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout gnd sky130_fd_pr__nfet_01v8 w=60 l=15
X2351 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2352 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2353 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 gnd sky130_fd_pr__res_generic_nd w=27 l=124
X2354 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 inp2 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2355 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2356 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2357 7bitdac_layout_1/x1_vref5 7bitdac_layout_1/x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
X2358 x1_vref5 x2_vref1 gnd sky130_fd_pr__res_generic_nd w=29 l=65
C0 d5 d4 20.96fF
C1 d6 d4 4.58fF
C2 d5 d6 10.80fF
C3 x1_out_v 7bitdac_layout_0/x1_out_v 2.44fF
C4 vdd d0 13.34fF
C5 vdd d1 10.67fF
C6 vdd d2 4.44fF
C7 7bitdac_layout_0/x1_out_v x2_vref1 12.72fF
C8 d1 d0 31.56fF
C9 d3 d1 6.49fF
C10 d2 d0 5.96fF
C11 d2 d1 17.88fF
C12 d3 d2 25.03fF
C13 d4 d3 21.63fF
C14 d4 d2 6.91fF
C15 d5 d0 2.75fF
C16 d6 d0 7.00fF
C17 d5 d3 5.61fF
C18 d6 d1 3.72fF
C19 vdd gnd 485.21fF
C20 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C21 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C22 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C23 7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C24 7bitdac_layout_1/x1_vref5 gnd 2.08fF
C25 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C26 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C27 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C28 7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C29 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C30 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C31 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C32 7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C33 7bitdac_layout_0/x1_vref5 gnd 2.08fF
C34 d0 gnd 228.24fF
C35 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C36 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C37 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 gnd 2.13fF
C38 7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 gnd 2.13fF
C39 d5 gnd 128.77fF
C40 d6 gnd 63.75fF
