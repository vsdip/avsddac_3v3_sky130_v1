magic
tech sky130A
magscale 1 2
timestamp 1640022418
<< error_p >>
rect 238 -246 280 -188
rect 528 -240 570 -184
<< ndiff >>
rect 238 -200 280 -188
rect 238 -234 242 -200
rect 276 -234 280 -200
rect 238 -246 280 -234
rect 528 -195 570 -184
rect 528 -229 532 -195
rect 566 -229 570 -195
rect 528 -240 570 -229
<< ndiffc >>
rect 242 -234 276 -200
rect 532 -229 566 -195
<< ndiffres >>
rect 228 -158 416 -156
rect 228 -184 596 -158
rect 228 -188 528 -184
rect 228 -246 238 -188
rect 280 -240 528 -188
rect 570 -240 596 -184
rect 280 -246 596 -240
rect 228 -284 596 -246
rect 416 -286 596 -284
<< locali >>
rect 224 -94 290 -90
rect 218 -200 308 -94
rect 218 -234 242 -200
rect 276 -234 308 -200
rect 218 -284 308 -234
rect 508 -195 598 -96
rect 508 -229 532 -195
rect 566 -229 598 -195
rect 508 -288 598 -229
<< end >>
