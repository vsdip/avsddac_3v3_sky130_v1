magic
tech sky130A
timestamp 1615764517
<< ndiffc >>
rect 119 -123 140 -94
rect 205 -124 226 -93
<< ndiffres >>
rect 114 -93 241 -78
rect 114 -94 205 -93
rect 114 -123 119 -94
rect 140 -123 205 -94
rect 114 -124 205 -123
rect 226 -124 241 -93
rect 114 -126 241 -124
rect 114 -142 242 -126
<< locali >>
rect 112 -47 145 -45
rect 109 -94 154 -47
rect 109 -123 119 -94
rect 140 -123 154 -94
rect 109 -142 154 -123
rect 195 -93 241 -77
rect 195 -124 205 -93
rect 226 -124 241 -93
rect 195 -171 241 -124
<< end >>
