magic
tech sky130A
timestamp 1616477680
<< locali >>
rect 151 11827 179 11867
rect 8205 6546 9704 6578
rect 9679 6525 9704 6546
rect 6872 6462 6931 6512
rect 6872 3296 6895 6462
rect 9679 6341 9706 6525
rect 9679 5974 9710 6341
rect 9679 5796 9712 5974
rect 9679 5599 9708 5796
rect 9679 5416 9710 5599
rect 9679 5034 9708 5416
rect 9679 4837 9706 5034
rect 9679 4665 9712 4837
rect 9679 4473 9708 4665
rect 9679 3519 9706 4473
rect 9683 3332 9710 3519
rect 6864 3289 6905 3296
rect 6864 3269 6875 3289
rect 6896 3269 6905 3289
rect 6864 3261 6905 3269
rect 5376 3088 5529 3159
rect 6869 3099 6910 3104
rect 5376 3086 5466 3088
rect 5376 2424 5422 3086
rect 6869 3074 6876 3099
rect 6900 3074 6910 3099
rect 6869 3069 6910 3074
rect 5385 2402 5422 2424
rect 5385 2011 5424 2402
rect 5385 1990 5401 2011
rect 5421 1990 5424 2011
rect 5385 1973 5424 1990
rect 3664 1702 3734 1743
rect 3665 1636 3730 1702
rect 5388 1658 5427 1687
rect 5388 1637 5392 1658
rect 5412 1637 5427 1658
rect 3663 1151 3732 1636
rect 3663 1130 3687 1151
rect 3704 1130 3732 1151
rect 3663 1113 3732 1130
rect 5388 1502 5427 1637
rect 1931 631 1968 886
rect 5388 781 5424 1502
rect 1931 609 1941 631
rect 1959 609 1968 631
rect 1931 597 1968 609
rect 3674 727 3732 772
rect 3674 706 3694 727
rect 3711 706 3732 727
rect 403 267 432 452
rect 403 247 409 267
rect 429 247 432 267
rect 403 243 432 247
rect 1931 402 1973 414
rect 1931 380 1940 402
rect 1958 380 1973 402
rect 403 166 432 171
rect 403 144 406 166
rect 427 144 432 166
rect 5 -56 40 10
rect -122 -90 40 -56
rect 5 -91 40 -90
rect 403 -87 432 144
rect 403 -104 408 -87
rect 426 -104 432 -87
rect 403 -108 432 -104
rect -35 -225 129 -193
rect 1931 -216 1973 380
rect 402 -247 431 -233
rect 402 -264 408 -247
rect 426 -264 431 -247
rect 1931 -238 1946 -216
rect 1964 -238 1973 -216
rect 1931 -264 1973 -238
rect 3674 -139 3732 706
rect 5388 348 5427 781
rect 5388 -7 5428 348
rect 5387 -28 5428 -7
rect 402 -519 431 -264
rect 1931 -475 1973 -458
rect 1931 -497 1941 -475
rect 1959 -497 1973 -475
rect 1931 -779 1973 -497
rect 3674 -520 3743 -139
rect 3674 -541 3706 -520
rect 3723 -541 3743 -520
rect 3674 -560 3743 -541
rect 3684 -822 3743 -800
rect 3684 -843 3707 -822
rect 3724 -843 3743 -822
rect 3684 -1365 3743 -843
rect 5386 -1095 5428 -28
rect 5386 -1116 5396 -1095
rect 5416 -1116 5428 -1095
rect 5386 -1128 5428 -1116
rect 5390 -1374 5429 -1370
rect 5390 -1406 5432 -1374
rect 5390 -1427 5403 -1406
rect 5423 -1427 5432 -1406
rect 5390 -2887 5432 -1427
rect 6874 -2224 6897 3069
rect 9683 2768 9708 3332
rect 9683 2571 9706 2768
rect 9683 2382 9708 2571
rect 9683 2202 9710 2382
rect 9683 1678 9712 2202
rect 9683 1481 9706 1678
rect 9683 1122 9710 1481
rect 9683 940 9708 1122
rect 9683 594 9706 940
rect 9679 553 9706 594
rect 9679 397 9704 553
rect 9775 255 9858 259
rect 9775 234 9779 255
rect 9797 234 9858 255
rect 9775 228 9858 234
rect 8554 150 8595 196
rect 9711 -10 9766 21
rect 6876 -2350 6896 -2224
rect 6875 -2356 6896 -2350
rect 6875 -2497 6895 -2356
rect 6874 -2503 6895 -2497
rect 6874 -2765 6894 -2503
rect 6867 -2775 6906 -2765
rect 6867 -2794 6878 -2775
rect 6897 -2794 6906 -2775
rect 6867 -2807 6906 -2794
rect 5390 -2925 5444 -2887
rect 6865 -2900 6904 -2888
rect 6865 -2921 6878 -2900
rect 6896 -2921 6904 -2900
rect 6865 -2930 6904 -2921
rect 6874 -3098 6894 -2930
rect 6874 -3106 6896 -3098
rect 6875 -5513 6896 -3106
rect 9736 -5444 9766 -10
rect 8160 -5486 9766 -5444
rect 8160 -5487 9733 -5486
rect 6875 -5517 6914 -5513
rect 6875 -5559 6896 -5517
rect 6875 -5563 6909 -5559
rect -45 -12065 -16 -12007
<< viali >>
rect 6875 3269 6896 3289
rect 6876 3074 6900 3099
rect 5401 1990 5421 2011
rect 5392 1637 5412 1658
rect 3687 1130 3704 1151
rect 1941 609 1959 631
rect 3694 706 3711 727
rect 409 247 429 267
rect 1940 380 1958 402
rect 406 144 427 166
rect 408 -104 426 -87
rect 408 -264 426 -247
rect 1946 -238 1964 -216
rect 1941 -497 1959 -475
rect 3706 -541 3723 -520
rect 3707 -843 3724 -822
rect 5396 -1116 5416 -1095
rect 5403 -1427 5423 -1406
rect 9779 234 9797 255
rect 6878 -2794 6897 -2775
rect 6878 -2921 6896 -2900
<< metal1 >>
rect 6864 3289 6905 3296
rect 6864 3269 6875 3289
rect 6896 3269 6905 3289
rect 6864 3261 6905 3269
rect 6875 3104 6895 3261
rect 6869 3099 6910 3104
rect 6869 3074 6876 3099
rect 6900 3074 6910 3099
rect 6869 3069 6910 3074
rect 6875 3066 6895 3069
rect 5385 2011 5424 2049
rect 5385 1990 5401 2011
rect 5421 1990 5424 2011
rect 5385 1709 5424 1990
rect 5388 1703 5424 1709
rect 5388 1658 5427 1703
rect 5388 1637 5392 1658
rect 5412 1637 5427 1658
rect 5388 1513 5427 1637
rect 3663 1151 3732 1188
rect 3663 1130 3687 1151
rect 3704 1130 3732 1151
rect 3663 727 3732 1130
rect 3663 706 3694 727
rect 3711 706 3732 727
rect 3663 665 3732 706
rect 1931 631 1968 645
rect 1931 609 1941 631
rect 1959 609 1968 631
rect 1931 402 1968 609
rect 1931 380 1940 402
rect 1958 380 1968 402
rect 9005 417 9059 420
rect 9005 384 9019 417
rect 9049 384 9059 417
rect 9005 380 9059 384
rect 1931 356 1968 380
rect 402 267 434 277
rect 402 247 409 267
rect 429 247 434 267
rect 9795 255 9804 259
rect 402 245 434 247
rect 404 174 433 245
rect 9797 234 9804 255
rect 9795 231 9804 234
rect 403 166 433 174
rect 403 164 406 166
rect 402 144 406 164
rect 427 145 433 166
rect 427 144 430 145
rect 402 143 430 144
rect 403 133 430 143
rect 8626 24 8684 51
rect 8626 -9 8638 24
rect 8669 -9 8684 24
rect 8626 -20 8684 -9
rect 402 -87 433 -80
rect 402 -95 408 -87
rect 403 -104 408 -95
rect 426 -95 433 -87
rect 426 -104 432 -95
rect 403 -247 432 -104
rect 403 -264 408 -247
rect 426 -264 432 -247
rect 403 -277 432 -264
rect 1931 -216 1973 -193
rect 1931 -238 1946 -216
rect 1964 -238 1973 -216
rect 1931 -475 1973 -238
rect 1931 -497 1941 -475
rect 1959 -497 1973 -475
rect 1931 -514 1973 -497
rect 3679 -520 3748 -475
rect 3679 -541 3706 -520
rect 3723 -541 3748 -520
rect 3679 -822 3748 -541
rect 3679 -843 3707 -822
rect 3724 -843 3748 -822
rect 3679 -896 3748 -843
rect 5386 -1095 5433 -1058
rect 5386 -1116 5396 -1095
rect 5416 -1116 5433 -1095
rect 5386 -1134 5433 -1116
rect 5385 -1329 5433 -1134
rect 5385 -1374 5429 -1329
rect 5385 -1406 5432 -1374
rect 5385 -1427 5403 -1406
rect 5423 -1427 5432 -1406
rect 5385 -1456 5432 -1427
rect 6867 -2775 6906 -2765
rect 6867 -2794 6878 -2775
rect 6897 -2794 6906 -2775
rect 6867 -2807 6906 -2794
rect 6874 -2888 6894 -2807
rect 6865 -2900 6904 -2888
rect 6865 -2921 6878 -2900
rect 6896 -2921 6904 -2900
rect 6865 -2930 6904 -2921
<< via1 >>
rect 9019 384 9049 417
rect 8638 -9 8669 24
<< metal2 >>
rect 6724 2529 8397 2582
rect 8343 25 8393 2529
rect 9014 458 9060 470
rect 9014 451 9024 458
rect 9015 425 9024 451
rect 9054 425 9060 458
rect 9015 417 9060 425
rect 9015 384 9019 417
rect 9049 384 9060 417
rect 9015 380 9060 384
rect 8636 25 8677 26
rect 8343 24 8677 25
rect 8343 0 8638 24
rect 8343 -2172 8393 0
rect 8636 -9 8638 0
rect 8669 -9 8677 24
rect 8636 -14 8677 -9
rect 8340 -3429 8397 -2172
rect 8340 -3486 8404 -3429
rect 8343 -3667 8404 -3486
rect 6685 -3720 8404 -3667
rect 8343 -3734 8404 -3720
<< via2 >>
rect 9024 425 9054 458
<< metal3 >>
rect 9015 525 9060 531
rect 9015 485 9022 525
rect 9055 485 9060 525
rect 9015 458 9060 485
rect 9015 425 9024 458
rect 9054 425 9060 458
rect 9015 422 9060 425
<< via3 >>
rect 9022 485 9055 525
<< metal4 >>
rect 8720 3561 9056 3562
rect 8295 3560 9056 3561
rect 7945 3558 9056 3560
rect 7561 3557 9056 3558
rect 6734 3553 9056 3557
rect 6325 3550 9056 3553
rect 5921 3526 9056 3550
rect 5921 3525 8390 3526
rect 5921 3523 8006 3525
rect 5921 3522 7586 3523
rect 5921 3518 6770 3522
rect 5921 3515 6366 3518
rect 9015 1734 9056 3526
rect 9015 1699 9058 1734
rect 9015 1270 9062 1699
rect 9016 1078 9062 1270
rect 8986 1075 9062 1078
rect 7334 1049 9062 1075
rect 7330 1035 9062 1049
rect 7330 -4617 7383 1035
rect 8986 1034 9062 1035
rect 9016 911 9062 1034
rect 9015 903 9062 911
rect 9015 538 9061 903
rect 9015 525 9060 538
rect 9015 485 9022 525
rect 9055 485 9060 525
rect 9015 481 9060 485
rect 7330 -4652 7392 -4617
rect 7334 -5130 7392 -4652
use 5bitdac_layout  5bitdac_layout_1
timestamp 1616476746
transform 1 0 -16 0 1 -5989
box -35 -6035 8186 5886
use 5bitdac_layout  5bitdac_layout_0
timestamp 1616476746
transform 1 0 34 0 1 6035
box -35 -6035 8186 5886
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 8567 0 1 -111
box 20 86 1230 590
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 -231 0 1 -33
box 109 -171 242 -45
<< labels >>
rlabel locali 9833 247 9833 247 1 out_v
rlabel locali 8569 165 8569 165 1 d5
rlabel locali 9692 524 9692 524 1 x1_out_v
rlabel locali 9757 -63 9757 -63 1 x2_out_v
rlabel locali -80 -76 -80 -76 1 x1_vref5
rlabel locali 32 -214 32 -214 1 x2_vref1
rlabel locali -33 -12045 -33 -12045 1 inp2
rlabel locali 161 11856 161 11856 1 inp1
rlabel locali 417 29 417 29 1 d0
rlabel locali 1956 -29 1956 -29 1 d1
rlabel locali 3703 -29 3703 -29 1 d2
rlabel locali 5399 -309 5399 -309 1 d3
rlabel locali 6883 -367 6883 -367 1 d4
rlabel metal4 9034 625 9034 625 1 vdd!
rlabel metal2 8370 10 8370 10 1 gnd!
<< end >>
