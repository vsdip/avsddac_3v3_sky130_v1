magic
tech sky130A
timestamp 1624221218
<< checkpaint >>
rect -521 -801 872 585
<< ndiff >>
rect 119 -100 140 -94
rect 119 -117 121 -100
rect 138 -117 140 -100
rect 119 -123 140 -117
rect 205 -100 226 -93
rect 205 -117 207 -100
rect 224 -117 226 -100
rect 205 -124 226 -117
<< ndiffc >>
rect 121 -117 138 -100
rect 207 -117 224 -100
<< ndiffres >>
rect 114 -93 241 -78
rect 114 -94 205 -93
rect 114 -123 119 -94
rect 140 -123 205 -94
rect 114 -124 205 -123
rect 226 -124 241 -93
rect 114 -126 241 -124
rect 114 -142 242 -126
<< locali >>
rect 112 -47 145 -45
rect 109 -100 154 -47
rect 109 -117 121 -100
rect 138 -117 154 -100
rect 109 -142 154 -117
rect 195 -100 241 -77
rect 195 -117 207 -100
rect 224 -117 241 -100
rect 195 -171 241 -117
<< end >>
