magic
tech sky130A
timestamp 1615766096
<< ndiffc >>
rect 119 -123 140 -94
rect 264 -120 285 -92
<< ndiffres >>
rect 114 -79 208 -78
rect 114 -92 298 -79
rect 114 -94 264 -92
rect 114 -123 119 -94
rect 140 -120 264 -94
rect 285 -120 298 -92
rect 140 -123 298 -120
rect 114 -142 298 -123
rect 208 -143 298 -142
<< locali >>
rect 112 -47 145 -45
rect 109 -94 154 -47
rect 109 -123 119 -94
rect 140 -123 154 -94
rect 109 -142 154 -123
rect 254 -92 299 -48
rect 254 -120 264 -92
rect 285 -120 299 -92
rect 254 -144 299 -120
<< end >>
