magic
tech sky130A
timestamp 1616555653
<< locali >>
rect 71802 26378 86734 26379
rect 71802 26359 99205 26378
rect 60161 26357 99205 26359
rect 60161 26337 71824 26357
rect 86727 26356 99205 26357
rect 48559 26291 48634 26292
rect 60161 26291 60182 26337
rect 48559 26289 60182 26291
rect 48559 26270 48565 26289
rect 48587 26270 60182 26289
rect 48559 26265 60182 26270
rect 48559 26264 60180 26265
rect 48140 26231 48171 26233
rect 49358 26231 49441 26233
rect 35727 26227 42825 26228
rect 47429 26227 48056 26228
rect 34699 26225 48056 26227
rect 34201 26224 48056 26225
rect 33828 26223 33855 26224
rect 34201 26223 48026 26224
rect 33828 26217 48026 26223
rect 33828 26200 33831 26217
rect 33848 26205 48026 26217
rect 48048 26205 48056 26224
rect 48129 26227 49441 26231
rect 48129 26208 48140 26227
rect 48162 26208 49441 26227
rect 48129 26207 49441 26208
rect 48129 26206 48756 26207
rect 33848 26204 48056 26205
rect 33848 26203 35732 26204
rect 42811 26203 48056 26204
rect 33848 26201 34723 26203
rect 48020 26201 48054 26203
rect 48140 26202 48171 26206
rect 33848 26200 34225 26201
rect 33828 26199 34225 26200
rect 33828 26196 33855 26199
rect 48559 26162 48592 26167
rect 48559 26143 48565 26162
rect 48587 26143 48592 26162
rect 398 25946 427 25977
rect 33825 25832 33855 25837
rect 33825 25815 33832 25832
rect 33849 25815 33855 25832
rect 33825 25808 33855 25815
rect 33829 23767 33850 25808
rect 33829 20919 33851 23767
rect 33829 20903 33852 20919
rect 33830 18070 33852 20903
rect 33829 18055 33852 18070
rect 33829 12378 33851 18055
rect 48559 14666 48592 26143
rect 49410 26124 49439 26207
rect 49411 25873 49439 26124
rect 48556 14143 48592 14666
rect 99180 14652 99205 26356
rect 99180 14645 99206 14652
rect 99181 14314 99206 14645
rect 48247 14108 48592 14143
rect 99180 14296 99206 14314
rect 46872 14044 46997 14068
rect 46874 13788 46915 14044
rect 95937 14007 96000 14014
rect 95937 13959 96004 14007
rect 95938 13957 95992 13959
rect 46874 13766 46886 13788
rect 46907 13766 46915 13788
rect 46874 13752 46915 13766
rect 95940 13924 95971 13957
rect 95940 13703 95969 13924
rect 95940 13684 95945 13703
rect 95963 13684 95969 13703
rect 95940 13680 95969 13684
rect 97257 13640 97274 14070
rect 99180 13855 99205 14296
rect 99264 13722 99305 13723
rect 99263 13716 99386 13722
rect 99263 13693 99268 13716
rect 99291 13693 99386 13716
rect 99263 13690 99386 13693
rect 99264 13687 99305 13690
rect 46874 13595 46917 13605
rect 46874 13573 46885 13595
rect 46906 13573 46917 13595
rect 46874 13244 46917 13573
rect 96050 13525 96076 13528
rect 95940 13519 96076 13525
rect 95940 13501 95946 13519
rect 95963 13501 96076 13519
rect 97257 13506 97276 13640
rect 98049 13609 98095 13655
rect 95940 13496 96076 13501
rect 46876 13218 46915 13244
rect 46874 13142 46915 13218
rect 33829 12366 33852 12378
rect 33830 9523 33852 12366
rect 33829 8373 33852 9523
rect 33829 8360 33853 8373
rect 33830 7224 33853 8360
rect 33830 6525 33854 7224
rect 33829 6514 33854 6525
rect 33829 5827 33853 6514
rect 33829 5815 33854 5827
rect 33830 3725 33854 5815
rect 33829 3715 33854 3725
rect 33829 3021 33853 3715
rect 33828 3015 33853 3021
rect 33828 2317 33852 3015
rect 33827 2311 33852 2317
rect 33827 1615 33851 2311
rect 33931 1752 34015 1764
rect 33930 1745 34015 1752
rect 33930 1643 33954 1745
rect 33827 1471 33852 1615
rect 34016 1471 34042 1545
rect 33827 1447 34042 1471
rect 33827 1445 34041 1447
rect 46874 1226 46900 13142
rect 82995 1633 83024 1686
rect 46871 1214 46900 1226
rect 34375 45 34408 50
rect 34375 20 34379 45
rect 34402 20 34408 45
rect 34375 15 34408 20
rect 34375 14 34409 15
rect 34380 9 34409 14
rect 34381 -113 34409 9
rect 34381 -926 34404 -113
rect 34379 -960 34404 -926
rect 35902 -915 35925 106
rect 37647 -857 37685 207
rect 39286 -810 39312 289
rect 40854 -751 40889 392
rect 42553 -645 42584 484
rect 45184 226 45220 589
rect 45180 172 45220 226
rect 45180 -521 45219 172
rect 46871 -434 46893 1214
rect 56387 938 56419 992
rect 56388 933 56419 938
rect 56388 916 56395 933
rect 56412 930 56419 933
rect 56412 916 56420 930
rect 56388 913 56420 916
rect 56388 912 56419 913
rect 52834 732 52877 750
rect 52834 708 52841 732
rect 52866 708 52877 732
rect 52834 698 52877 708
rect 96050 599 96076 13496
rect 97253 13399 97278 13506
rect 97253 13397 97983 13399
rect 99190 13397 99215 13480
rect 97253 13370 99215 13397
rect 97253 13366 99211 13370
rect 97780 13364 99211 13366
rect 49669 116 49703 568
rect 52829 504 52869 516
rect 54575 509 54600 510
rect 51188 484 51227 503
rect 51188 464 51199 484
rect 51221 464 51227 484
rect 52829 480 52836 504
rect 52861 480 52869 504
rect 52829 476 52869 480
rect 54574 504 54600 509
rect 54574 486 54578 504
rect 54596 486 54600 504
rect 54574 480 54600 486
rect 56390 484 56419 498
rect 51188 236 51227 464
rect 49669 -380 49701 116
rect 51188 -321 51222 236
rect 52835 67 52857 476
rect 51188 -341 51193 -321
rect 51215 -341 51222 -321
rect 51188 -357 51222 -341
rect 52836 -375 52857 67
rect 54574 -342 54598 480
rect 56390 467 56397 484
rect 56414 467 56419 484
rect 56390 114 56419 467
rect 57817 453 57867 464
rect 57817 428 57830 453
rect 57854 428 57867 453
rect 57817 229 57867 428
rect 56388 29 56419 114
rect 57814 137 57867 229
rect 56388 -330 56417 29
rect 49669 -401 49673 -380
rect 49692 -401 49701 -380
rect 49669 -404 49701 -401
rect 52835 -381 52870 -375
rect 52835 -402 52839 -381
rect 52861 -402 52870 -381
rect 54574 -380 54600 -342
rect 56388 -347 56396 -330
rect 56413 -347 56417 -330
rect 57814 -346 57864 137
rect 56388 -355 56417 -347
rect 57813 -358 57864 -346
rect 57813 -365 57831 -358
rect 54574 -397 54577 -380
rect 54596 -397 54600 -380
rect 57814 -383 57831 -365
rect 57855 -383 57864 -358
rect 57814 -388 57864 -383
rect 54574 -400 54600 -397
rect 52835 -407 52870 -402
rect 96045 -415 96081 599
rect 96045 -430 96079 -415
rect 94389 -434 96079 -430
rect 46871 -454 96079 -434
rect 45180 -548 70599 -521
rect 45180 -567 70565 -548
rect 70584 -567 70599 -548
rect 45180 -584 70599 -567
rect 45180 -589 45219 -584
rect 42552 -648 47892 -645
rect 42552 -650 53233 -648
rect 42552 -652 56617 -650
rect 42552 -658 57864 -652
rect 42552 -679 57826 -658
rect 42553 -680 42584 -679
rect 47865 -682 57826 -679
rect 53216 -683 57826 -682
rect 57850 -683 57864 -658
rect 53216 -688 57864 -683
rect 56604 -692 57864 -688
rect 40856 -761 40889 -751
rect 40856 -764 43555 -761
rect 46224 -764 56416 -761
rect 40856 -766 56416 -764
rect 40856 -783 56397 -766
rect 56414 -783 56416 -766
rect 40856 -789 56416 -783
rect 43540 -792 46246 -789
rect 39286 -811 39377 -810
rect 40873 -811 40901 -808
rect 45344 -811 47373 -810
rect 54575 -811 54605 -806
rect 39285 -828 54578 -811
rect 54597 -828 54605 -811
rect 39285 -829 54605 -828
rect 39285 -830 45355 -829
rect 54573 -834 54605 -829
rect 37762 -857 52861 -855
rect 37647 -862 52861 -857
rect 37647 -875 52834 -862
rect 37647 -876 39311 -875
rect 37647 -883 37879 -876
rect 52827 -886 52834 -875
rect 52856 -886 52861 -862
rect 52827 -891 52861 -886
rect 52827 -894 52858 -891
rect 37831 -909 51042 -907
rect 35902 -916 35999 -915
rect 37831 -916 51216 -909
rect 35902 -918 51216 -916
rect 35902 -938 51190 -918
rect 51212 -938 51216 -918
rect 35902 -939 51216 -938
rect 35973 -941 51216 -939
rect 37831 -943 51216 -941
rect 51027 -945 51216 -943
rect 34379 -961 49695 -960
rect 34379 -978 49671 -961
rect 34380 -981 49671 -978
rect 35972 -982 49671 -981
rect 49690 -982 49695 -961
rect 35972 -983 49695 -982
rect 49665 -988 49694 -983
<< viali >>
rect 48565 26270 48587 26289
rect 33831 26200 33848 26217
rect 48026 26205 48048 26224
rect 48140 26208 48162 26227
rect 48565 26143 48587 26162
rect 33832 25815 33849 25832
rect 46886 13766 46907 13788
rect 95945 13684 95963 13703
rect 99268 13693 99291 13716
rect 46885 13573 46906 13595
rect 95946 13501 95963 13519
rect 34379 20 34402 45
rect 57830 1198 57854 1223
rect 56395 916 56412 933
rect 54579 835 54597 853
rect 52841 708 52866 732
rect 51199 597 51221 617
rect 51199 464 51221 484
rect 52836 480 52861 504
rect 54578 486 54596 504
rect 51193 -341 51215 -321
rect 56397 467 56414 484
rect 70569 466 70588 485
rect 57830 428 57854 453
rect 49673 -401 49692 -380
rect 52839 -402 52861 -381
rect 56396 -347 56413 -330
rect 54577 -397 54596 -380
rect 57831 -383 57855 -358
rect 70565 -567 70584 -548
rect 57826 -683 57850 -658
rect 56397 -783 56414 -766
rect 54578 -828 54597 -811
rect 52834 -886 52856 -862
rect 51190 -938 51212 -918
rect 49671 -982 49690 -961
<< metal1 >>
rect 48559 26289 48593 26293
rect 48559 26270 48565 26289
rect 48587 26270 48593 26289
rect 48559 26264 48593 26270
rect 48140 26231 48171 26233
rect 48019 26227 48171 26231
rect 48019 26224 48140 26227
rect 33828 26217 33855 26224
rect 33828 26200 33831 26217
rect 33848 26200 33855 26217
rect 48019 26205 48026 26224
rect 48048 26208 48140 26224
rect 48162 26208 48171 26227
rect 48048 26205 48171 26208
rect 48019 26203 48171 26205
rect 48020 26201 48054 26203
rect 48140 26202 48171 26203
rect 33828 26196 33855 26200
rect 33829 25837 33850 26196
rect 48559 26164 48592 26264
rect 48559 26162 48593 26164
rect 48559 26143 48565 26162
rect 48587 26143 48593 26162
rect 48559 26135 48593 26143
rect 33825 25832 33855 25837
rect 33825 25815 33832 25832
rect 33849 25815 33855 25832
rect 33825 25808 33855 25815
rect 98503 13870 98558 13874
rect 98503 13844 98522 13870
rect 98550 13844 98558 13870
rect 98503 13840 98558 13844
rect 46875 13788 46917 13799
rect 46875 13766 46886 13788
rect 46907 13766 46917 13788
rect 46875 13595 46917 13766
rect 99264 13716 99305 13723
rect 46875 13573 46885 13595
rect 46906 13573 46917 13595
rect 46875 13566 46917 13573
rect 95940 13703 95969 13709
rect 95940 13684 95945 13703
rect 95963 13684 95969 13703
rect 99264 13693 99268 13716
rect 99291 13693 99305 13716
rect 99264 13687 99305 13693
rect 95940 13680 95969 13684
rect 95940 13525 95968 13680
rect 95940 13519 95969 13525
rect 95940 13501 95946 13519
rect 95963 13501 95969 13519
rect 95940 13496 95969 13501
rect 98141 13486 98186 13512
rect 98141 13453 98147 13486
rect 98177 13453 98186 13486
rect 98141 13443 98186 13453
rect 57817 1223 57861 1253
rect 57817 1198 57830 1223
rect 57854 1198 57861 1223
rect 56388 935 56419 937
rect 56388 933 56420 935
rect 56388 916 56395 933
rect 56412 916 56420 933
rect 56388 913 56420 916
rect 54575 853 54600 862
rect 54575 835 54579 853
rect 54597 835 54600 853
rect 52834 732 52877 750
rect 52834 708 52841 732
rect 52866 708 52877 732
rect 52834 698 52877 708
rect 34374 50 34408 656
rect 51191 617 51232 630
rect 51191 597 51199 617
rect 51221 597 51232 617
rect 51191 484 51232 597
rect 52834 516 52855 698
rect 51191 464 51199 484
rect 51221 464 51232 484
rect 52829 504 52869 516
rect 54575 509 54600 835
rect 52829 480 52836 504
rect 52861 480 52869 504
rect 54574 504 54600 509
rect 54574 486 54578 504
rect 54596 486 54600 504
rect 54574 480 54600 486
rect 56388 484 56417 913
rect 52829 476 52869 480
rect 51191 448 51232 464
rect 56388 467 56397 484
rect 56414 467 56417 484
rect 56388 460 56417 467
rect 57817 453 57861 1198
rect 57817 428 57830 453
rect 57854 428 57861 453
rect 57817 414 57861 428
rect 70551 485 70602 587
rect 70551 466 70569 485
rect 70588 466 70602 485
rect 34375 45 34408 50
rect 34375 20 34379 45
rect 34402 20 34408 45
rect 34375 14 34408 20
rect 51185 -321 51219 -303
rect 51185 -341 51193 -321
rect 51215 -341 51219 -321
rect 49664 -380 49696 -366
rect 49664 -401 49673 -380
rect 49692 -401 49696 -380
rect 49664 -952 49696 -401
rect 51185 -918 51219 -341
rect 56390 -330 56419 -315
rect 56390 -347 56396 -330
rect 56413 -347 56419 -330
rect 52835 -381 52870 -375
rect 52835 -402 52839 -381
rect 52861 -402 52870 -381
rect 52835 -407 52870 -402
rect 54574 -380 54600 -373
rect 54574 -397 54577 -380
rect 54596 -397 54600 -380
rect 54574 -400 54600 -397
rect 52836 -857 52857 -407
rect 54574 -806 54598 -400
rect 56390 -766 56419 -347
rect 57813 -358 57863 -346
rect 57813 -362 57831 -358
rect 57811 -383 57831 -362
rect 57855 -365 57863 -358
rect 57855 -383 57861 -365
rect 57811 -658 57861 -383
rect 70551 -515 70602 466
rect 70551 -548 70599 -515
rect 70551 -567 70565 -548
rect 70584 -567 70599 -548
rect 70551 -582 70599 -567
rect 57811 -683 57826 -658
rect 57850 -683 57861 -658
rect 57811 -689 57861 -683
rect 56390 -783 56397 -766
rect 56414 -783 56419 -766
rect 56390 -790 56419 -783
rect 54574 -811 54605 -806
rect 54574 -820 54578 -811
rect 54573 -828 54578 -820
rect 54597 -828 54605 -811
rect 54573 -834 54605 -828
rect 52830 -860 52861 -857
rect 52827 -862 52861 -860
rect 52827 -886 52834 -862
rect 52856 -886 52861 -862
rect 52827 -891 52861 -886
rect 52827 -894 52858 -891
rect 51185 -938 51190 -918
rect 51212 -938 51219 -918
rect 51185 -945 51219 -938
rect 49664 -961 49695 -952
rect 49664 -973 49671 -961
rect 49665 -982 49671 -973
rect 49690 -982 49695 -961
rect 49665 -983 49695 -982
rect 49665 -988 49694 -983
<< via1 >>
rect 98522 13844 98550 13870
rect 98147 13453 98177 13486
<< metal2 >>
rect 54482 25959 54543 25965
rect 54479 25941 54543 25959
rect 39303 25870 39868 25872
rect 54479 25871 54508 25941
rect 50304 25870 54508 25871
rect 39303 25850 54508 25870
rect 39303 25847 54500 25850
rect 39306 22792 39333 25847
rect 98515 13912 98560 13913
rect 98515 13881 98524 13912
rect 98554 13881 98560 13912
rect 98515 13870 98560 13881
rect 98515 13844 98522 13870
rect 98550 13844 98560 13870
rect 98515 13840 98560 13844
rect 95969 13665 97424 13667
rect 95969 13644 97908 13665
rect 97407 13643 97908 13644
rect 97877 13481 97908 13643
rect 98099 13486 98181 13492
rect 98099 13481 98147 13486
rect 97877 13453 98147 13481
rect 98177 13453 98181 13486
rect 97877 13443 98181 13453
rect 97877 13435 98116 13443
<< via2 >>
rect 98524 13881 98554 13912
<< metal3 >>
rect 98515 13959 98560 13970
rect 98515 13924 98522 13959
rect 98559 13924 98560 13959
rect 98515 13913 98560 13924
rect 98516 13912 98560 13913
rect 98516 13881 98524 13912
rect 98554 13881 98560 13912
rect 98516 13878 98560 13881
<< via3 >>
rect 98522 13924 98559 13959
<< metal4 >>
rect 49359 25879 50242 25914
rect 49360 25747 49403 25879
rect 49362 25698 49400 25747
rect 50198 25702 50238 25879
rect 38239 25602 41487 25603
rect 49362 25602 49398 25698
rect 38239 25567 49398 25602
rect 96420 14615 96634 14616
rect 98349 14615 98568 14621
rect 96420 14580 98570 14615
rect 98349 14578 98570 14580
rect 98522 13990 98570 14578
rect 98516 13979 98570 13990
rect 98516 13959 98564 13979
rect 98516 13924 98522 13959
rect 98559 13924 98564 13959
rect 98516 13917 98564 13924
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 33821 0 1 1698
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 98066 0 1 13350
box 20 86 1230 590
use 8bitdac_layout  8bitdac_layout_1
timestamp 1616493856
transform 1 0 49013 0 1 543
box 0 -616 48260 25781
use 8bitdac_layout  8bitdac_layout_0
timestamp 1616493856
transform 1 0 0 0 1 616
box 0 -616 48260 25781
<< labels >>
rlabel locali 99333 13702 99333 13702 1 out_v
rlabel metal4 98536 13979 98536 13979 1 vdd!
rlabel metal2 98121 13464 98121 13464 1 gnd!
rlabel locali 99198 13397 99198 13397 1 x2_out_v
rlabel locali 99196 13952 99196 13952 1 x1_out_v
rlabel locali 98070 13633 98070 13633 1 d8
rlabel locali 33943 1696 33943 1696 1 x1_vref5
rlabel locali 34028 1477 34028 1477 1 x2_vref1
rlabel locali 83006 1654 83006 1654 1 inp2
rlabel locali 412 25966 412 25966 1 inp1
rlabel locali 34390 -33 34390 -33 1 d0
rlabel locali 45207 291 45207 291 1 d6
rlabel locali 46882 1330 46882 1330 1 d7
rlabel locali 42567 -454 42567 -454 1 d5
rlabel locali 40873 -670 40873 -670 1 d4
rlabel locali 39297 -242 39297 -242 1 d3
rlabel locali 37666 -769 37666 -769 1 d2
rlabel locali 35912 -810 35912 -810 1 d1
<< end >>
