magic
tech sky130A
timestamp 1616567895
<< viali >>
rect 102718 28781 102738 28799
<< metal1 >>
rect 102715 28807 102801 28812
rect 102715 28799 102773 28807
rect 102715 28781 102718 28799
rect 102738 28781 102773 28799
rect 102715 28779 102773 28781
rect 102800 28779 102801 28807
rect 102715 28774 102801 28779
rect 104169 26312 104281 26348
<< via1 >>
rect 102773 28779 102800 28807
<< metal2 >>
rect 102769 28810 102861 28813
rect 102769 28807 102824 28810
rect 102769 28779 102773 28807
rect 102800 28779 102824 28807
rect 102769 28778 102824 28779
rect 102855 28778 102861 28810
rect 102769 28774 102861 28778
<< via2 >>
rect 102824 28778 102855 28810
<< metal3 >>
rect 102875 28816 102931 28819
rect 102819 28814 102931 28816
rect 102819 28810 102884 28814
rect 102819 28778 102824 28810
rect 102855 28778 102884 28810
rect 102919 28778 102931 28814
rect 102819 28774 102931 28778
rect 102875 28773 102931 28774
rect 104169 26312 104281 26348
<< via3 >>
rect 102884 28778 102919 28814
<< mimcapcontact >>
rect 105103 28779 105138 28813
<< metal4 >>
rect 102882 28814 105143 28816
rect 102882 28778 102884 28814
rect 102919 28813 105143 28814
rect 102919 28779 105103 28813
rect 105138 28779 105143 28813
rect 102919 28778 105143 28779
rect 102882 28776 105143 28778
rect 102882 28774 102978 28776
use cap_28p  cap_28p_0
timestamp 1616448691
transform 1 0 105249 0 1 26963
box -984 -1226 12410 12449
use 10bitdac_layout  10bitdac_layout_0
timestamp 1616566027
transform 1 0 214 0 1 28846
box -214 -28846 102528 27385
<< labels >>
rlabel metal3 104180 26326 104180 26326 1 gnd!
rlabel metal4 103604 28795 103604 28795 1 out_v
<< end >>
