magic
tech sky130A
timestamp 1615739263
<< nwell >>
rect 253 311 301 586
rect 583 327 774 550
rect 908 86 1100 312
<< nmos >>
rect 1005 410 1020 470
rect 675 170 690 230
<< pmos >>
rect 675 350 690 471
rect 1005 165 1020 285
<< ndiff >>
rect 960 456 1005 470
rect 960 425 965 456
rect 990 425 1005 456
rect 960 410 1005 425
rect 1020 456 1065 470
rect 1020 425 1035 456
rect 1060 425 1065 456
rect 1020 410 1065 425
rect 630 215 675 230
rect 630 185 635 215
rect 659 185 675 215
rect 630 170 675 185
rect 690 216 735 230
rect 690 184 705 216
rect 730 184 735 216
rect 690 170 735 184
<< pdiff >>
rect 635 438 675 471
rect 635 379 640 438
rect 660 379 675 438
rect 635 350 675 379
rect 690 440 731 471
rect 690 380 705 440
rect 725 380 731 440
rect 690 350 731 380
rect 965 254 1005 285
rect 965 194 970 254
rect 990 194 1005 254
rect 965 165 1005 194
rect 1020 255 1061 285
rect 1020 195 1035 255
rect 1055 195 1061 255
rect 1020 165 1061 195
<< ndiffc >>
rect 965 425 990 456
rect 1035 425 1060 456
rect 635 185 659 215
rect 705 184 730 216
<< pdiffc >>
rect 640 379 660 438
rect 705 380 725 440
rect 970 194 990 254
rect 1035 195 1055 255
<< poly >>
rect 675 471 690 485
rect 1005 470 1020 485
rect 1005 395 1020 410
rect 1085 409 1115 420
rect 1085 395 1091 409
rect 1004 389 1091 395
rect 1109 389 1115 409
rect 1004 380 1115 389
rect 460 290 492 291
rect 365 280 492 290
rect 365 271 467 280
rect 460 260 467 271
rect 485 260 492 280
rect 460 252 492 260
rect 595 288 624 291
rect 675 288 690 350
rect 595 280 690 288
rect 1005 285 1020 380
rect 595 260 600 280
rect 618 270 690 280
rect 618 260 624 270
rect 595 252 624 260
rect 675 230 690 270
rect 675 155 690 170
rect 1005 149 1020 165
<< polycont >>
rect 1091 389 1109 409
rect 467 260 485 280
rect 600 260 618 280
<< locali >>
rect 246 496 306 571
rect 615 505 1140 535
rect 635 438 660 505
rect 635 379 640 438
rect 635 350 660 379
rect 705 440 731 472
rect 725 380 731 440
rect 421 340 422 341
rect 420 335 435 340
rect 395 315 405 324
rect 425 315 435 335
rect 20 259 98 306
rect 395 305 417 315
rect 420 311 435 315
rect 705 311 731 380
rect 960 456 990 470
rect 960 425 965 456
rect 960 365 990 425
rect 1035 456 1065 505
rect 1060 425 1065 456
rect 1035 410 1065 425
rect 1085 415 1115 420
rect 1085 409 1175 415
rect 1085 389 1091 409
rect 1109 407 1175 409
rect 1109 389 1152 407
rect 1169 389 1175 407
rect 1085 380 1175 389
rect 704 305 731 311
rect 859 344 966 365
rect 983 344 990 365
rect 859 339 990 344
rect 859 305 890 339
rect 207 271 285 290
rect 460 280 624 291
rect 460 260 467 280
rect 485 260 600 280
rect 618 260 624 280
rect 704 276 890 305
rect 704 275 735 276
rect 859 275 890 276
rect 460 252 624 260
rect 630 215 660 230
rect 630 185 635 215
rect 659 185 660 215
rect 251 96 311 156
rect 630 130 660 185
rect 705 216 735 275
rect 730 184 735 216
rect 705 170 735 184
rect 965 254 990 339
rect 965 194 970 254
rect 965 165 990 194
rect 1035 255 1061 285
rect 1055 195 1061 255
rect 1035 130 1061 195
rect 625 100 1150 130
<< viali >>
rect 405 315 425 335
rect 1152 389 1169 407
rect 966 344 983 365
<< metal1 >>
rect 251 490 301 575
rect 519 574 1165 590
rect 519 569 1166 574
rect 520 460 540 569
rect 460 440 540 460
rect 460 340 480 440
rect 1146 415 1166 569
rect 1146 407 1175 415
rect 1146 389 1152 407
rect 1169 389 1175 407
rect 1146 385 1175 389
rect 960 365 1230 370
rect 960 344 966 365
rect 983 344 1230 365
rect 960 340 1230 344
rect 395 335 480 340
rect 395 315 405 335
rect 425 315 480 335
rect 395 311 480 315
rect 256 91 306 162
use INV  INV_1
timestamp 1615514756
transform 1 0 301 0 1 311
box -44 -220 145 275
use INV  INV_0
timestamp 1615514756
transform 1 0 112 0 1 311
box -44 -220 145 275
<< labels >>
rlabel metal1 272 534 272 534 1 vdd!
rlabel metal1 270 108 270 108 1 gnd!
rlabel locali 788 110 788 110 1 inp2
rlabel locali 889 516 889 516 1 inp1
rlabel locali 50 283 50 283 1 din
rlabel space 373 298 373 298 1 dinb
rlabel locali 235 278 235 278 1 dinb
rlabel space 413 298 413 298 1 dd
rlabel poly 1058 388 1058 388 1 dd
rlabel metal1 1056 351 1056 351 1 vout
<< end >>
