magic
tech sky130A
magscale 1 2
timestamp 1625518311
<< locali >>
rect 46054 508408 47990 508612
rect 1388 508124 18224 508148
rect 1040 508082 18224 508124
rect 34048 508082 47990 508408
rect 1040 508050 47990 508082
rect 1040 508016 1076 508050
rect 1110 508016 47990 508050
rect 1040 507948 47990 508016
rect 1388 507936 47990 507948
rect 17790 507870 47990 507936
rect 34048 507680 47990 507870
rect 41820 465164 42396 465210
rect 12010 464980 36218 465044
rect 41796 464980 42534 465164
rect 1308 464958 1904 464962
rect 12010 464958 42534 464980
rect 1308 464938 42534 464958
rect 1280 464892 42534 464938
rect 1280 464786 1317 464892
rect 1423 464786 42534 464892
rect 1280 464720 42534 464786
rect 1308 464718 42534 464720
rect 1308 464714 12998 464718
rect 1734 464688 12998 464714
rect 35038 464634 42534 464718
rect 41796 464282 42534 464634
rect 41820 464174 42454 464282
rect 41936 442502 42454 464174
rect 46054 443352 47990 507680
rect 41950 426232 42396 442502
rect 46152 426512 47038 443352
rect 41660 426014 42778 426232
rect 41660 425188 41849 426014
rect 42675 425188 42778 426014
rect 41660 424942 42778 425188
rect 45470 425825 48130 426512
rect 41950 424874 42396 424942
rect 45470 423919 45929 425825
rect 47547 423919 48130 425825
rect 45470 423444 48130 423919
rect 86114 421766 86752 421910
rect 40164 421718 44794 421764
rect 47536 421718 87094 421766
rect 31504 421694 87094 421718
rect 12258 421678 87094 421694
rect 1326 421674 87094 421678
rect 1052 421608 87094 421674
rect 1052 421574 1082 421608
rect 1116 421574 87094 421608
rect 1052 421516 87094 421574
rect 1326 421510 87094 421516
rect 1326 421494 31986 421510
rect 12258 421486 31986 421494
rect 40164 421482 44794 421510
rect 47536 421488 87094 421510
rect 86080 420832 86752 421488
rect 41660 419072 42846 419336
rect 41660 418390 41899 419072
rect 42581 418390 42846 419072
rect 41660 418178 42846 418390
rect 41942 416032 42480 418178
rect 35606 378752 36994 378954
rect 14172 378540 36994 378752
rect 1396 378492 1600 378500
rect 1786 378492 36994 378540
rect 1396 378402 36994 378492
rect 1396 378368 1451 378402
rect 1485 378368 36994 378402
rect 1396 378264 36994 378368
rect 1786 378236 36994 378264
rect 14172 378112 36994 378236
rect 32172 335486 32496 335558
rect 28860 335424 32496 335486
rect 10856 335392 32496 335424
rect 1434 335252 1730 335338
rect 6558 335272 32496 335392
rect 2098 335252 32496 335272
rect 1434 335240 32496 335252
rect 1434 335062 1470 335240
rect 1648 335174 32496 335240
rect 1648 335074 7088 335174
rect 10856 335112 29920 335174
rect 1648 335062 1730 335074
rect 1434 334992 1730 335062
rect 2098 335054 7088 335074
rect 32172 334974 32496 335174
rect 32172 322958 32560 334974
rect 32106 322634 32560 322958
rect 32106 294014 32236 322634
rect 32106 292560 32348 294014
rect 28540 292024 28614 292088
rect 28256 292012 28622 292024
rect 1210 292006 1346 292008
rect 1708 292006 28622 292012
rect 1210 291982 28622 292006
rect 1210 291948 1250 291982
rect 1284 291948 28622 291982
rect 1210 291910 28622 291948
rect 1210 291876 1250 291910
rect 1284 291876 28622 291910
rect 1210 291848 28622 291876
rect 1238 291840 28622 291848
rect 1708 291776 28622 291840
rect 1708 291750 28614 291776
rect 28500 291716 28614 291750
rect 1478 248988 2134 248998
rect 1478 248986 2176 248988
rect 1478 248946 13250 248986
rect 27000 248976 27368 249020
rect 27000 248964 27428 248976
rect 20984 248962 27428 248964
rect 20984 248946 27057 248962
rect 1478 248917 27057 248946
rect 1478 248883 1504 248917
rect 1538 248883 1576 248917
rect 1610 248883 27057 248917
rect 1478 248822 27057 248883
rect 1478 248820 2176 248822
rect 1520 248810 2176 248820
rect 12604 248784 27057 248822
rect 27307 248784 27428 248962
rect 12604 248782 27428 248784
rect 27000 248722 27428 248782
rect 27000 248690 27368 248722
rect 28540 235124 28614 291716
rect 32122 265398 32348 292560
rect 32122 264580 32380 265398
rect 32154 250476 32380 264580
rect 32090 250284 32380 250476
rect 29152 248914 29456 248964
rect 29152 248736 29220 248914
rect 29398 248736 29456 248914
rect 29152 248706 29456 248736
rect 28540 235100 28634 235124
rect 28580 234270 28634 235100
rect 29192 234566 29314 248706
rect 32090 235686 32316 250284
rect 35606 249642 36994 378112
rect 41950 366394 42396 416032
rect 45196 414571 47856 415122
rect 45196 412665 45757 414571
rect 47375 412665 47856 414571
rect 45196 412054 47856 412665
rect 45264 386360 45606 412054
rect 41894 366122 42396 366394
rect 45196 384980 45606 386360
rect 41894 289002 42340 366122
rect 45196 295526 45600 384980
rect 86080 306970 86664 420832
rect 86080 303878 86746 306970
rect 45154 295098 45600 295526
rect 42024 256962 42302 289002
rect 35376 249272 36994 249642
rect 41996 256738 42302 256962
rect 35376 235714 36648 249272
rect 41996 245398 42274 256738
rect 45154 250810 45558 295098
rect 86366 284952 86746 303878
rect 86330 284286 86746 284952
rect 86330 262694 86710 284286
rect 86266 262268 86710 262694
rect 45154 249138 45752 250810
rect 41968 244896 42274 245398
rect 41968 236116 42246 244896
rect 41940 235758 42246 236116
rect 32090 235362 32418 235686
rect 29174 234444 29314 234566
rect 32152 234446 32418 235362
rect 35676 234936 36022 235714
rect 41940 235030 42230 235758
rect 45248 235474 45752 249138
rect 86266 240392 86646 262268
rect 86266 240010 86738 240392
rect 86418 235878 86738 240010
rect 86388 235814 86738 235878
rect 86388 235638 86676 235814
rect 45250 235167 45618 235474
rect 86388 235460 86463 235638
rect 86569 235460 86676 235638
rect 86388 235434 86676 235460
rect 45250 235061 45339 235167
rect 45517 235061 45618 235167
rect 35678 234648 35914 234936
rect 41940 234861 42236 235030
rect 45250 235016 45618 235061
rect 45250 234948 45614 235016
rect 41940 234755 42024 234861
rect 42130 234755 42236 234861
rect 41940 234676 42236 234755
rect 35654 234583 35986 234648
rect 35654 234477 35717 234583
rect 35895 234477 35986 234583
rect 29174 234216 29266 234444
rect 32152 234430 32434 234446
rect 32156 234369 32434 234430
rect 35654 234422 35986 234477
rect 32156 234263 32246 234369
rect 32352 234263 32434 234369
rect 29158 234188 29278 234216
rect 29158 234154 29199 234188
rect 29233 234154 29278 234188
rect 32156 234174 32434 234263
rect 29158 234124 29278 234154
rect 41944 233739 42200 233802
rect 29162 233686 29262 233712
rect 29162 233652 29196 233686
rect 29230 233652 29262 233686
rect 29162 233630 29262 233652
rect 41944 233633 42006 233739
rect 42112 233633 42200 233739
rect 29184 233074 29246 233630
rect 41944 233564 42200 233633
rect 45254 233655 45620 233742
rect 32254 233244 32334 233256
rect 32220 233191 32390 233244
rect 32220 233157 32250 233191
rect 32284 233157 32322 233191
rect 32356 233157 32390 233191
rect 32220 233116 32390 233157
rect 28944 232638 28982 232674
rect 32254 232594 32334 233116
rect 35696 232627 35934 232672
rect 28750 232528 28856 232566
rect 28750 232494 28785 232528
rect 28819 232494 28856 232528
rect 28750 232468 28856 232494
rect 35696 232521 35765 232627
rect 35871 232521 35934 232627
rect 35696 232470 35934 232521
rect 35756 231476 35846 232470
rect 41998 228770 42132 233564
rect 45254 233477 45343 233655
rect 45521 233477 45620 233655
rect 86392 233741 86686 233800
rect 86392 233635 86457 233741
rect 86563 233635 86686 233741
rect 86392 233562 86686 233635
rect 45254 233422 45620 233477
rect 41992 228688 42160 228770
rect 41992 228654 42046 228688
rect 42080 228654 42160 228688
rect 41992 228598 42160 228654
rect 45314 228638 45568 233422
rect 86446 232544 86604 233562
rect 86436 232032 86632 232544
rect 86436 231926 86484 232032
rect 86590 231926 86632 232032
rect 86436 231880 86632 231926
rect 86428 228906 86626 228948
rect 86428 228800 86475 228906
rect 86581 228800 86626 228906
rect 86428 228756 86626 228800
rect 41990 228340 42160 228376
rect 41990 228306 42048 228340
rect 42082 228306 42160 228340
rect 41990 228234 42160 228306
rect 42036 223014 42082 228234
rect 45318 223760 45474 228638
rect 86474 228184 86574 228756
rect 45240 223688 45566 223760
rect 45240 223582 45302 223688
rect 45480 223582 45566 223688
rect 45240 223512 45566 223582
rect 45318 223014 45474 223022
rect 45260 222954 45534 223014
rect 45260 222848 45330 222954
rect 45436 222848 45534 222954
rect 45260 222790 45534 222848
rect 45318 217796 45474 222790
rect 45308 217598 45474 217796
rect 45308 212510 45464 217598
rect 45306 212372 45464 212510
rect 45306 210400 45426 212372
rect 45306 210354 45466 210400
rect 45412 210352 45466 210354
rect 230072 179868 230166 180094
rect 230074 179422 230156 179868
rect 230074 179324 230166 179422
rect 230082 177260 230166 179324
rect 230084 176058 230162 177260
rect 230080 173642 230200 176058
rect 230046 158416 230234 173642
rect 230036 158212 230234 158416
rect 230036 152361 230218 158212
rect 230036 152255 230079 152361
rect 230185 152255 230218 152361
rect 230036 152248 230218 152255
rect 230040 152206 230212 152248
rect 223454 151670 223526 151896
rect 223390 151658 223526 151670
rect 223390 151624 223403 151658
rect 223437 151624 223526 151658
rect 223390 151618 223526 151624
rect 230050 151745 230232 151788
rect 230050 151639 230087 151745
rect 230193 151639 230232 151745
rect 223394 151218 223516 151236
rect 223394 151184 223405 151218
rect 223439 151184 223516 151218
rect 223394 151168 223516 151184
rect 223464 151058 223516 151168
rect 230050 151124 230232 151639
rect 223464 150824 223514 151058
rect 223466 150572 223508 150824
rect 223464 150556 223508 150572
rect 223464 150150 223506 150556
rect 223464 144986 223528 150150
rect 223464 141836 223524 144986
rect 215750 123988 215830 125568
rect 215722 123944 215860 123988
rect 215722 123910 215774 123944
rect 215808 123910 215860 123944
rect 215722 123854 215860 123910
rect 215750 123852 215830 123854
rect 215722 123506 215860 123558
rect 215722 123472 215770 123506
rect 215804 123472 215860 123506
rect 215722 123424 215860 123472
rect 215744 122952 215830 123424
rect 219388 123230 219598 123902
rect 215644 121622 215932 122952
rect 157096 121566 200074 121594
rect 213632 121566 216026 121622
rect 34792 121478 39042 121506
rect 45868 121478 50118 121536
rect 157096 121478 216026 121566
rect 13216 121448 17466 121478
rect 34792 121448 50118 121478
rect 61214 121448 65464 121478
rect 68830 121448 73080 121478
rect 94098 121448 98348 121478
rect 101712 121448 113520 121478
rect 153316 121448 216026 121478
rect 5658 121424 17466 121448
rect 1760 121420 17466 121424
rect 24264 121420 28514 121448
rect 31504 121420 73080 121448
rect 90262 121420 113520 121448
rect 116338 121420 123876 121448
rect 1760 121414 73080 121420
rect 1326 121392 73080 121414
rect 75608 121392 83146 121420
rect 86166 121392 123876 121420
rect 126894 121392 131144 121448
rect 138288 121420 146288 121448
rect 149510 121420 216026 121448
rect 138288 121392 216026 121420
rect 1326 121299 216026 121392
rect 1326 121265 1377 121299
rect 1411 121276 216026 121299
rect 1411 121265 35754 121276
rect 1326 121248 35754 121265
rect 38312 121248 216026 121276
rect 1326 121218 13572 121248
rect 17052 121218 35754 121248
rect 46474 121218 62148 121248
rect 65166 121218 69416 121248
rect 71714 121218 102126 121248
rect 112760 121218 153760 121248
rect 157096 121218 216026 121248
rect 1326 121194 6010 121218
rect 1326 121192 1940 121194
rect 17052 121190 24850 121218
rect 27898 121190 32148 121218
rect 46474 121190 50724 121218
rect 71714 121190 90416 121218
rect 71714 121162 75964 121190
rect 82762 121162 87012 121190
rect 94126 121132 98376 121218
rect 112760 121190 117010 121218
rect 123462 121162 127712 121218
rect 130702 121162 138674 121218
rect 145760 121190 150010 121218
rect 199556 121190 216026 121218
rect 219390 115908 219452 123230
rect 219376 110454 219472 115908
rect 219376 110292 219554 110454
rect 219384 82632 219554 110292
rect 1322 78178 2024 78182
rect 1322 78162 2042 78178
rect 1322 78120 7396 78162
rect 107308 78120 108944 78276
rect 219344 78120 219688 82632
rect 1322 78094 108944 78120
rect 1322 78060 1379 78094
rect 1413 78060 108944 78094
rect 1322 78022 108944 78060
rect 1322 77988 1379 78022
rect 1413 77988 108944 78022
rect 1322 77946 108944 77988
rect 1340 77944 108944 77946
rect 1340 77942 3194 77944
rect 1792 77924 3194 77942
rect 6570 77912 108944 77944
rect 107308 77846 108944 77912
rect 205854 77846 220472 78120
rect 107068 77638 220472 77846
rect 107308 77500 108944 77638
rect 205854 77316 220472 77638
rect 219344 77296 219688 77316
rect 223440 52746 223570 141836
rect 230044 91166 230250 151124
rect 25162 34966 135052 34980
rect 1442 34914 2048 34926
rect 2804 34914 135052 34966
rect 1442 34842 135052 34914
rect 1442 34808 1473 34842
rect 1507 34808 135052 34842
rect 1442 34754 135052 34808
rect 223418 34774 223602 52746
rect 1442 34736 2934 34754
rect 1442 34732 2048 34736
rect 25162 34696 135052 34754
rect 222918 34696 223756 34774
rect 133346 34554 223756 34696
rect 222918 34460 223756 34554
rect 223418 34408 223602 34460
rect 230038 24152 230352 91166
rect 10676 13808 11714 13994
rect 230054 13866 230334 24152
rect 229026 13808 230364 13866
rect 10676 13562 230364 13808
rect 2508 13548 230364 13562
rect 1320 13494 230364 13548
rect 1048 13429 230364 13494
rect 1048 13395 1073 13429
rect 1107 13395 230364 13429
rect 1048 13336 230364 13395
rect 1054 13334 230364 13336
rect 1320 13322 230364 13334
rect 2508 13310 230364 13322
rect 2508 13292 12146 13310
rect 10676 13016 11714 13292
rect 229026 13274 230364 13310
rect 230054 13182 230334 13274
<< viali >>
rect 1076 508016 1110 508050
rect 1317 464786 1423 464892
rect 41849 425188 42675 426014
rect 45929 423919 47547 425825
rect 1082 421574 1116 421608
rect 41899 418390 42581 419072
rect 1451 378368 1485 378402
rect 1470 335062 1648 335240
rect 1250 291948 1284 291982
rect 1250 291876 1284 291910
rect 1504 248883 1538 248917
rect 1576 248883 1610 248917
rect 27057 248784 27307 248962
rect 29220 248736 29398 248914
rect 45757 412665 47375 414571
rect 86463 235460 86569 235638
rect 45339 235061 45517 235167
rect 42024 234755 42130 234861
rect 35717 234477 35895 234583
rect 32246 234263 32352 234369
rect 29199 234154 29233 234188
rect 29196 233652 29230 233686
rect 42006 233633 42112 233739
rect 32250 233157 32284 233191
rect 32322 233157 32356 233191
rect 28785 232494 28819 232528
rect 35765 232521 35871 232627
rect 45343 233477 45521 233655
rect 86457 233635 86563 233741
rect 42046 228654 42080 228688
rect 86484 231926 86590 232032
rect 86475 228800 86581 228906
rect 42048 228306 42082 228340
rect 45302 223582 45480 223688
rect 45330 222848 45436 222954
rect 230079 152255 230185 152361
rect 223403 151624 223437 151658
rect 230087 151639 230193 151745
rect 223405 151184 223439 151218
rect 215774 123910 215808 123944
rect 215770 123472 215804 123506
rect 1377 121265 1411 121299
rect 1379 78060 1413 78094
rect 1379 77988 1413 78022
rect 1473 34808 1507 34842
rect 1073 13395 1107 13429
<< metal1 >>
rect 674 508061 1152 508092
rect 674 508009 691 508061
rect 743 508009 755 508061
rect 807 508050 1152 508061
rect 807 508016 1076 508050
rect 1110 508016 1152 508050
rect 807 508009 1152 508016
rect 674 507972 1152 508009
rect 858 464901 1446 464918
rect 858 464785 880 464901
rect 996 464892 1446 464901
rect 996 464786 1317 464892
rect 1423 464786 1446 464892
rect 996 464785 1446 464786
rect 858 464744 1446 464785
rect 41688 426014 42818 426226
rect 41688 425188 41849 426014
rect 42675 425188 42818 426014
rect 744 421621 1154 421646
rect 744 421569 776 421621
rect 828 421608 1154 421621
rect 828 421574 1082 421608
rect 1116 421574 1154 421608
rect 828 421569 1154 421574
rect 744 421538 1154 421569
rect 41688 419072 42818 425188
rect 45402 425825 48130 426308
rect 45402 424738 45929 425825
rect 41688 418390 41899 419072
rect 42581 418390 42818 419072
rect 41688 418094 42818 418390
rect 45264 423919 45929 424738
rect 47547 423919 48130 425825
rect 45264 423512 48130 423919
rect 45264 415122 47514 423512
rect 45196 414571 47856 415122
rect 45196 412665 45757 414571
rect 47375 412665 47856 414571
rect 45196 412054 47856 412665
rect 1372 378452 1536 378454
rect 812 378404 1536 378452
rect 812 378352 849 378404
rect 901 378352 913 378404
rect 965 378402 1536 378404
rect 965 378368 1451 378402
rect 1485 378368 1536 378402
rect 965 378352 1536 378368
rect 812 378310 1536 378352
rect 736 335276 980 335306
rect 736 335240 1676 335276
rect 736 335210 1470 335240
rect 736 335094 800 335210
rect 916 335094 1470 335210
rect 736 335062 1470 335094
rect 1648 335062 1676 335240
rect 736 335030 1676 335062
rect 736 335014 980 335030
rect 832 291997 1318 292004
rect 832 291945 863 291997
rect 915 291982 1318 291997
rect 915 291948 1250 291982
rect 1284 291948 1318 291982
rect 915 291945 1318 291948
rect 832 291933 1318 291945
rect 832 291881 863 291933
rect 915 291910 1318 291933
rect 915 291881 1250 291910
rect 832 291876 1250 291881
rect 1284 291876 1318 291910
rect 832 291854 1318 291876
rect 840 248936 1632 248964
rect 840 248884 856 248936
rect 908 248884 920 248936
rect 972 248917 1632 248936
rect 972 248884 1504 248917
rect 840 248883 1504 248884
rect 1538 248883 1576 248917
rect 1610 248883 1632 248917
rect 840 248840 1632 248883
rect 26962 248962 29600 249046
rect 26962 248784 27057 248962
rect 27307 248914 29600 248962
rect 27307 248784 29220 248914
rect 26962 248736 29220 248784
rect 29398 248736 29600 248914
rect 26962 248618 29600 248736
rect 86404 235638 86644 235662
rect 86404 235460 86463 235638
rect 86569 235460 86644 235638
rect 86404 235360 86644 235460
rect 86402 235332 86644 235360
rect 45264 235167 45628 235248
rect 45264 235061 45339 235167
rect 45517 235061 45628 235167
rect 41960 234861 42190 234940
rect 41960 234755 42024 234861
rect 42130 234755 42190 234861
rect 45264 234796 45628 235061
rect 35682 234583 35936 234634
rect 35682 234477 35717 234583
rect 35895 234477 35936 234583
rect 32196 234369 32414 234418
rect 32196 234263 32246 234369
rect 32352 234263 32414 234369
rect 35682 234324 35936 234477
rect 29148 234188 29288 234220
rect 29148 234154 29199 234188
rect 29233 234154 29288 234188
rect 29148 234128 29288 234154
rect 29146 234104 29288 234128
rect 32196 234206 32414 234263
rect 35678 234260 35936 234324
rect 41960 234620 42190 234755
rect 29146 233686 29276 234104
rect 32196 234102 32406 234206
rect 29146 233652 29196 233686
rect 29230 233652 29276 233686
rect 29146 233622 29276 233652
rect 32212 233256 32390 234102
rect 32204 233191 32398 233256
rect 32204 233157 32250 233191
rect 32284 233157 32322 233191
rect 32356 233157 32398 233191
rect 32204 233096 32398 233157
rect 35678 232627 35934 234260
rect 41960 233739 42186 234620
rect 45260 233742 45636 234796
rect 41960 233633 42006 233739
rect 42112 233633 42186 233739
rect 41960 233582 42186 233633
rect 45254 233655 45636 233742
rect 45254 233477 45343 233655
rect 45521 233498 45636 233655
rect 86402 233741 86638 235332
rect 86402 233635 86457 233741
rect 86563 233635 86638 233741
rect 86402 233570 86638 233635
rect 45521 233477 45620 233498
rect 45254 233422 45620 233477
rect 28750 232528 28862 232580
rect 28750 232494 28785 232528
rect 28819 232494 28862 232528
rect 28750 232466 28862 232494
rect 35678 232521 35765 232627
rect 35871 232521 35934 232627
rect 35678 232484 35934 232521
rect 28754 232194 28858 232466
rect 28744 232154 28882 232194
rect 28744 232102 28784 232154
rect 28836 232102 28882 232154
rect 28744 232058 28882 232102
rect 86416 232032 86666 232072
rect 86416 231926 86484 232032
rect 86590 231926 86666 232032
rect 86416 231876 86666 231926
rect 86438 228940 86616 231876
rect 86434 228906 86624 228940
rect 86434 228800 86475 228906
rect 86581 228800 86624 228906
rect 42012 228688 42114 228736
rect 86434 228704 86624 228800
rect 42012 228654 42046 228688
rect 42080 228654 42114 228688
rect 42012 228340 42114 228654
rect 42012 228306 42048 228340
rect 42082 228306 42114 228340
rect 42012 228260 42114 228306
rect 45254 223688 45552 223756
rect 45254 223582 45302 223688
rect 45480 223582 45552 223688
rect 45254 222954 45552 223582
rect 45254 222854 45330 222954
rect 45266 222848 45330 222854
rect 45436 222854 45552 222954
rect 45436 222848 45538 222854
rect 45266 222812 45538 222848
rect 230008 152361 230260 152390
rect 230008 152255 230079 152361
rect 230185 152255 230260 152361
rect 230008 151810 230260 152255
rect 230008 151745 230278 151810
rect 230008 151718 230087 151745
rect 223388 151658 223452 151670
rect 223388 151624 223403 151658
rect 223437 151624 223452 151658
rect 223388 151618 223452 151624
rect 230012 151639 230087 151718
rect 230193 151639 230278 151745
rect 223392 151236 223444 151618
rect 230012 151600 230278 151639
rect 223392 151218 223450 151236
rect 223392 151186 223405 151218
rect 223396 151184 223405 151186
rect 223439 151184 223450 151218
rect 223396 151168 223450 151184
rect 215720 123944 215896 123990
rect 215720 123910 215774 123944
rect 215808 123910 215896 123944
rect 215720 123506 215896 123910
rect 215720 123472 215770 123506
rect 215804 123472 215896 123506
rect 215720 123408 215896 123472
rect 730 121313 1458 121352
rect 730 121261 762 121313
rect 814 121261 826 121313
rect 878 121299 1458 121313
rect 878 121265 1377 121299
rect 1411 121265 1458 121299
rect 878 121261 1458 121265
rect 730 121218 1458 121261
rect 784 78094 1460 78116
rect 784 78067 1379 78094
rect 784 78015 796 78067
rect 848 78015 860 78067
rect 912 78060 1379 78067
rect 1413 78060 1460 78094
rect 912 78022 1460 78060
rect 912 78015 1379 78022
rect 784 77988 1379 78015
rect 1413 77988 1460 78022
rect 784 77972 1460 77988
rect 808 34859 1536 34878
rect 808 34807 849 34859
rect 901 34842 1536 34859
rect 901 34808 1473 34842
rect 1507 34808 1536 34842
rect 901 34807 1536 34808
rect 808 34770 1536 34807
rect 660 13438 1130 13460
rect 660 13386 702 13438
rect 754 13429 1130 13438
rect 754 13395 1073 13429
rect 1107 13395 1130 13429
rect 754 13386 1130 13395
rect 660 13360 1130 13386
<< via1 >>
rect 691 508009 743 508061
rect 755 508009 807 508061
rect 880 464785 996 464901
rect 776 421569 828 421621
rect 849 378352 901 378404
rect 913 378352 965 378404
rect 800 335094 916 335210
rect 863 291945 915 291997
rect 863 291881 915 291933
rect 856 248884 908 248936
rect 920 248884 972 248936
rect 28784 232102 28836 232154
rect 762 121261 814 121313
rect 826 121261 878 121313
rect 796 78015 848 78067
rect 860 78015 912 78067
rect 849 34807 901 34859
rect 702 13386 754 13438
<< metal2 >>
rect 342 508066 830 508114
rect 342 508010 376 508066
rect 432 508061 830 508066
rect 432 508010 691 508061
rect 342 508009 691 508010
rect 743 508009 755 508061
rect 807 508009 830 508061
rect 342 507944 830 508009
rect 796 464926 1006 464934
rect 326 464901 1006 464926
rect 326 464843 880 464901
rect 326 464787 377 464843
rect 433 464787 880 464843
rect 326 464785 880 464787
rect 996 464785 1006 464901
rect 326 464718 1006 464785
rect 374 421625 856 421668
rect 374 421569 396 421625
rect 452 421621 856 421625
rect 452 421569 776 421621
rect 828 421569 856 421621
rect 374 421522 856 421569
rect 308 378404 1008 378486
rect 308 378402 849 378404
rect 308 378346 378 378402
rect 434 378352 849 378402
rect 901 378352 913 378404
rect 965 378352 1008 378404
rect 434 378346 1008 378352
rect 308 378272 1008 378346
rect 296 335256 494 335298
rect 296 335210 968 335256
rect 296 335177 800 335210
rect 296 335121 369 335177
rect 425 335121 800 335177
rect 296 335094 800 335121
rect 916 335094 968 335210
rect 296 335058 968 335094
rect 296 335038 494 335058
rect 698 292000 938 292006
rect 320 291997 938 292000
rect 320 291963 863 291997
rect 320 291907 365 291963
rect 421 291945 863 291963
rect 915 291945 938 291997
rect 421 291933 938 291945
rect 421 291907 863 291933
rect 320 291881 863 291907
rect 915 291881 938 291933
rect 320 291862 938 291881
rect 302 248936 996 249006
rect 302 248934 856 248936
rect 302 248878 327 248934
rect 383 248878 407 248934
rect 463 248884 856 248934
rect 908 248884 920 248936
rect 972 248884 996 248936
rect 463 248878 996 248884
rect 302 248810 996 248878
rect 28748 232162 28880 232186
rect 28748 232154 29326 232162
rect 28748 232102 28784 232154
rect 28836 232102 29326 232154
rect 28748 232100 29326 232102
rect 28748 232096 28888 232100
rect 28748 232058 28880 232096
rect 2946 175569 4258 175780
rect 2946 174953 3108 175569
rect 3964 174953 4258 175569
rect 2946 174794 4258 174953
rect 2946 174760 7564 174794
rect 2946 174724 13834 174760
rect 2946 174700 21328 174724
rect 22726 174704 27330 174712
rect 22726 174700 28900 174704
rect 2946 174648 28900 174700
rect 2946 174636 22896 174648
rect 27278 174640 28900 174648
rect 2946 174620 13834 174636
rect 2946 174588 4258 174620
rect 7402 174588 13834 174620
rect 312 121313 898 121392
rect 312 121312 762 121313
rect 312 121256 365 121312
rect 421 121261 762 121312
rect 814 121261 826 121313
rect 878 121261 898 121313
rect 421 121256 898 121261
rect 312 121188 898 121256
rect 336 78089 924 78158
rect 336 78033 384 78089
rect 440 78067 924 78089
rect 440 78033 796 78067
rect 336 78015 796 78033
rect 848 78015 860 78067
rect 912 78015 924 78067
rect 336 77948 924 78015
rect 332 34869 954 34918
rect 332 34813 373 34869
rect 429 34859 954 34869
rect 429 34813 849 34859
rect 332 34807 849 34813
rect 901 34807 954 34859
rect 332 34744 954 34807
rect 328 13440 788 13494
rect 328 13384 370 13440
rect 426 13438 788 13440
rect 426 13386 702 13438
rect 754 13386 788 13438
rect 426 13384 788 13386
rect 328 13334 788 13384
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 376 508010 432 508066
rect 377 464787 433 464843
rect 396 421569 452 421625
rect 378 378346 434 378402
rect 369 335121 425 335177
rect 365 291907 421 291963
rect 327 248878 383 248934
rect 407 248878 463 248934
rect 3108 174953 3964 175569
rect 365 121256 421 121312
rect 384 78033 440 78089
rect 373 34813 429 34869
rect 370 13384 426 13440
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect -800 680242 1700 685242
rect 120410 679704 124992 702300
rect 120240 679290 124992 679704
rect 120240 677386 120858 679290
rect 124122 677386 124992 679290
rect 582300 677984 584800 682984
rect 120240 677350 124992 677386
rect 120240 676552 124950 677350
rect -800 645284 1660 648642
rect -800 644260 163 645284
rect 1347 644762 1660 645284
rect 1347 644336 30974 644762
rect 1347 644260 1660 644336
rect -800 643842 1660 644260
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 508066 480 508096
rect -800 508010 376 508066
rect 432 508010 480 508066
rect -800 507984 480 508010
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464843 480 464874
rect -800 464787 377 464843
rect 433 464787 480 464843
rect -800 464762 480 464787
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421625 480 421652
rect -800 421569 396 421625
rect 452 421569 480 421625
rect -800 421540 480 421569
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378402 480 378430
rect -800 378346 378 378402
rect 434 378346 480 378402
rect -800 378318 480 378346
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect 122 336274 478 336278
rect -800 335177 480 335208
rect -800 335121 369 335177
rect 425 335121 480 335177
rect -800 335096 480 335121
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291963 480 291986
rect -800 291907 365 291963
rect 421 291907 480 291963
rect -800 291874 480 291907
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248934 480 248964
rect -800 248878 327 248934
rect 383 248878 407 248934
rect 463 248878 480 248934
rect -800 248852 480 248878
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect -800 175696 1660 177688
rect -800 175569 4126 175696
rect -800 174953 3108 175569
rect 3964 174953 4126 175569
rect -800 174836 4126 174953
rect -800 172888 1660 174836
rect 233894 172718 265130 202950
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121312 480 121342
rect -800 121256 365 121312
rect 421 121256 480 121312
rect -800 121230 480 121256
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78089 480 78120
rect -800 78033 384 78089
rect 440 78033 480 78089
rect -800 78008 480 78033
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34869 480 34898
rect -800 34813 373 34869
rect 429 34813 480 34869
rect -800 34786 480 34813
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13440 480 13476
rect -800 13384 370 13440
rect 426 13384 480 13440
rect -800 13364 480 13384
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 120858 677386 124122 679290
rect 163 644260 1347 645284
<< mimcap >>
rect 235850 174040 262698 201416
<< metal4 >>
rect 120366 679290 125496 680040
rect 120366 679074 120858 679290
rect 120198 677386 120858 679074
rect 124122 679074 125496 679290
rect 124122 679062 127430 679074
rect 197836 679062 234588 679164
rect 124122 677386 234588 679062
rect 120198 677308 234588 677386
rect 120366 677286 234588 677308
rect 120366 677218 200848 677286
rect 120366 676720 125496 677218
rect -854 645284 2056 645488
rect -854 644260 163 645284
rect 1347 644762 2056 645284
rect 30512 644762 30990 646010
rect 1347 644336 30990 644762
rect 1347 644260 2056 644336
rect -854 644034 2056 644260
rect 30512 552250 30990 644336
rect 233136 562822 234460 677286
rect 30536 234560 30826 552250
rect 233136 545444 235866 562822
rect 233218 545114 235866 545444
rect 234388 494250 234710 545114
rect 234364 493666 234710 494250
rect 234364 431964 234686 493666
rect 234364 428392 234734 431964
rect 234524 330316 234734 428392
rect 234524 328398 234736 330316
rect 234526 278386 234736 328398
rect 234526 277472 234746 278386
rect 30402 234282 31114 234560
rect 30854 233842 30954 234282
rect 234536 226754 234746 277472
rect 234536 225542 234778 226754
rect 234542 204802 234778 225542
rect 234580 192660 234660 204802
rect 234580 192270 234700 192660
rect 234612 188780 234700 192270
rect 234602 188632 234700 188780
rect 234602 180872 234690 188632
rect 234606 180162 234670 180872
use 10bitdac_cap_layout_design  10bitdac_cap_layout_design_0
timestamp 1625518311
transform 1 0 27354 0 1 122658
box 0 -48 235318 112414
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 8338 0 0 0 gpio_analog[0]
flabel metal3 s -800 381864 480 381976 0 FreeSans 8338 0 0 0 gpio_analog[10]
flabel metal3 s -800 338642 480 338754 0 FreeSans 8338 0 0 0 gpio_analog[11]
flabel metal3 s -800 295420 480 295532 0 FreeSans 8338 0 0 0 gpio_analog[12]
flabel metal3 s -800 252398 480 252510 0 FreeSans 8338 0 0 0 gpio_analog[13]
flabel metal3 s -800 124776 480 124888 0 FreeSans 8338 0 0 0 gpio_analog[14]
flabel metal3 s -800 81554 480 81666 0 FreeSans 8338 0 0 0 gpio_analog[15]
flabel metal3 s -800 38332 480 38444 0 FreeSans 8338 0 0 0 gpio_analog[16]
flabel metal3 s -800 16910 480 17022 0 FreeSans 8338 0 0 0 gpio_analog[17]
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 8338 0 0 0 gpio_analog[1]
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 8338 0 0 0 gpio_analog[2]
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 8338 0 0 0 gpio_analog[3]
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 8338 0 0 0 gpio_analog[4]
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 8338 0 0 0 gpio_analog[5]
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 8338 0 0 0 gpio_analog[6]
flabel metal3 s -800 511530 480 511642 0 FreeSans 8338 0 0 0 gpio_analog[7]
flabel metal3 s -800 468308 480 468420 0 FreeSans 8338 0 0 0 gpio_analog[8]
flabel metal3 s -800 425086 480 425198 0 FreeSans 8338 0 0 0 gpio_analog[9]
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 8338 0 0 0 gpio_noesd[0]
flabel metal3 s -800 380682 480 380794 0 FreeSans 8338 0 0 0 gpio_noesd[10]
flabel metal3 s -800 337460 480 337572 0 FreeSans 8338 0 0 0 gpio_noesd[11]
flabel metal3 s -800 294238 480 294350 0 FreeSans 8338 0 0 0 gpio_noesd[12]
flabel metal3 s -800 251216 480 251328 0 FreeSans 8338 0 0 0 gpio_noesd[13]
flabel metal3 s -800 123594 480 123706 0 FreeSans 8338 0 0 0 gpio_noesd[14]
flabel metal3 s -800 80372 480 80484 0 FreeSans 8338 0 0 0 gpio_noesd[15]
flabel metal3 s -800 37150 480 37262 0 FreeSans 8338 0 0 0 gpio_noesd[16]
flabel metal3 s -800 15728 480 15840 0 FreeSans 8338 0 0 0 gpio_noesd[17]
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 8338 0 0 0 gpio_noesd[1]
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 8338 0 0 0 gpio_noesd[2]
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 8338 0 0 0 gpio_noesd[3]
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 8338 0 0 0 gpio_noesd[4]
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 8338 0 0 0 gpio_noesd[5]
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 8338 0 0 0 gpio_noesd[6]
flabel metal3 s -800 510348 480 510460 0 FreeSans 8338 0 0 0 gpio_noesd[7]
flabel metal3 s -800 467126 480 467238 0 FreeSans 8338 0 0 0 gpio_noesd[8]
flabel metal3 s -800 423904 480 424016 0 FreeSans 8338 0 0 0 gpio_noesd[9]
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 8338 0 0 0 io_analog[0]
flabel metal3 s 0 680242 1700 685242 0 FreeSans 8338 0 0 0 io_analog[10]
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 14300 180 0 0 io_analog[1]
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 14300 180 0 0 io_analog[2]
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 14300 180 0 0 io_analog[3]
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 14300 180 0 0 io_analog[4]
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 14300 180 0 0 io_analog[5]
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 14300 180 0 0 io_analog[6]
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 14300 180 0 0 io_analog[7]
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 14300 180 0 0 io_analog[8]
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 14300 180 0 0 io_analog[9]
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 14300 180 0 0 io_analog[4]
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 14300 180 0 0 io_analog[5]
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 14300 180 0 0 io_analog[6]
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 14300 180 0 0 io_clamp_high[0]
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 14300 180 0 0 io_clamp_high[1]
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 14300 180 0 0 io_clamp_high[2]
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 14300 180 0 0 io_clamp_low[0]
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 14300 180 0 0 io_clamp_low[1]
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 14300 180 0 0 io_clamp_low[2]
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 8338 0 0 0 io_in[0]
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 8338 0 0 0 io_in[10]
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 8338 0 0 0 io_in[11]
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 8338 0 0 0 io_in[12]
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 8338 0 0 0 io_in[13]
flabel metal3 s -800 507984 480 508096 0 FreeSans 8338 0 0 0 io_in[14]
flabel metal3 s -800 464762 480 464874 0 FreeSans 8338 0 0 0 io_in[15]
flabel metal3 s -800 421540 480 421652 0 FreeSans 8338 0 0 0 io_in[16]
flabel metal3 s -800 378318 480 378430 0 FreeSans 8338 0 0 0 io_in[17]
flabel metal3 s -800 335096 480 335208 0 FreeSans 8338 0 0 0 io_in[18]
flabel metal3 s -800 291874 480 291986 0 FreeSans 8338 0 0 0 io_in[19]
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 8338 0 0 0 io_in[1]
flabel metal3 s -800 248852 480 248964 0 FreeSans 8338 0 0 0 io_in[20]
flabel metal3 s -800 121230 480 121342 0 FreeSans 8338 0 0 0 io_in[21]
flabel metal3 s -800 78008 480 78120 0 FreeSans 8338 0 0 0 io_in[22]
flabel metal3 s -800 34786 480 34898 0 FreeSans 8338 0 0 0 io_in[23]
flabel metal3 s -800 13364 480 13476 0 FreeSans 8338 0 0 0 io_in[24]
flabel metal3 s -800 8636 480 8748 0 FreeSans 8338 0 0 0 io_in[25]
flabel metal3 s -800 3908 480 4020 0 FreeSans 8338 0 0 0 io_in[26]
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 8338 0 0 0 io_in[2]
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 8338 0 0 0 io_in[3]
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 8338 0 0 0 io_in[4]
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 8338 0 0 0 io_in[5]
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 8338 0 0 0 io_in[6]
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 8338 0 0 0 io_in[7]
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 8338 0 0 0 io_in[8]
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 8338 0 0 0 io_in[9]
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 8338 0 0 0 io_in_3v3[0]
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 8338 0 0 0 io_in_3v3[10]
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 8338 0 0 0 io_in_3v3[11]
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 8338 0 0 0 io_in_3v3[12]
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 8338 0 0 0 io_in_3v3[13]
flabel metal3 s -800 509166 480 509278 0 FreeSans 8338 0 0 0 io_in_3v3[14]
flabel metal3 s -800 465944 480 466056 0 FreeSans 8338 0 0 0 io_in_3v3[15]
flabel metal3 s -800 422722 480 422834 0 FreeSans 8338 0 0 0 io_in_3v3[16]
flabel metal3 s -800 379500 480 379612 0 FreeSans 8338 0 0 0 io_in_3v3[17]
flabel metal3 s -800 336278 480 336390 0 FreeSans 8338 0 0 0 io_in_3v3[18]
flabel metal3 s -800 293056 480 293168 0 FreeSans 8338 0 0 0 io_in_3v3[19]
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 8338 0 0 0 io_in_3v3[1]
flabel metal3 s -800 250034 480 250146 0 FreeSans 8338 0 0 0 io_in_3v3[20]
flabel metal3 s -800 122412 480 122524 0 FreeSans 8338 0 0 0 io_in_3v3[21]
flabel metal3 s -800 79190 480 79302 0 FreeSans 8338 0 0 0 io_in_3v3[22]
flabel metal3 s -800 35968 480 36080 0 FreeSans 8338 0 0 0 io_in_3v3[23]
flabel metal3 s -800 14546 480 14658 0 FreeSans 8338 0 0 0 io_in_3v3[24]
flabel metal3 s -800 9818 480 9930 0 FreeSans 8338 0 0 0 io_in_3v3[25]
flabel metal3 s -800 5090 480 5202 0 FreeSans 8338 0 0 0 io_in_3v3[26]
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 8338 0 0 0 io_in_3v3[2]
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 8338 0 0 0 io_in_3v3[3]
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 8338 0 0 0 io_in_3v3[4]
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 8338 0 0 0 io_in_3v3[5]
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 8338 0 0 0 io_in_3v3[6]
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 8338 0 0 0 io_in_3v3[7]
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 8338 0 0 0 io_in_3v3[8]
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 8338 0 0 0 io_in_3v3[9]
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 8338 0 0 0 io_oeb[0]
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 8338 0 0 0 io_oeb[10]
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 8338 0 0 0 io_oeb[11]
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 8338 0 0 0 io_oeb[12]
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 8338 0 0 0 io_oeb[13]
flabel metal3 s -800 505620 480 505732 0 FreeSans 8338 0 0 0 io_oeb[14]
flabel metal3 s -800 462398 480 462510 0 FreeSans 8338 0 0 0 io_oeb[15]
flabel metal3 s -800 419176 480 419288 0 FreeSans 8338 0 0 0 io_oeb[16]
flabel metal3 s -800 375954 480 376066 0 FreeSans 8338 0 0 0 io_oeb[17]
flabel metal3 s -800 332732 480 332844 0 FreeSans 8338 0 0 0 io_oeb[18]
flabel metal3 s -800 289510 480 289622 0 FreeSans 8338 0 0 0 io_oeb[19]
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 8338 0 0 0 io_oeb[1]
flabel metal3 s -800 246488 480 246600 0 FreeSans 8338 0 0 0 io_oeb[20]
flabel metal3 s -800 118866 480 118978 0 FreeSans 8338 0 0 0 io_oeb[21]
flabel metal3 s -800 75644 480 75756 0 FreeSans 8338 0 0 0 io_oeb[22]
flabel metal3 s -800 32422 480 32534 0 FreeSans 8338 0 0 0 io_oeb[23]
flabel metal3 s -800 11000 480 11112 0 FreeSans 8338 0 0 0 io_oeb[24]
flabel metal3 s -800 6272 480 6384 0 FreeSans 8338 0 0 0 io_oeb[25]
flabel metal3 s -800 1544 480 1656 0 FreeSans 8338 0 0 0 io_oeb[26]
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 8338 0 0 0 io_oeb[2]
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 8338 0 0 0 io_oeb[3]
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 8338 0 0 0 io_oeb[4]
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 8338 0 0 0 io_oeb[5]
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 8338 0 0 0 io_oeb[6]
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 8338 0 0 0 io_oeb[7]
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 8338 0 0 0 io_oeb[8]
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 8338 0 0 0 io_oeb[9]
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 8338 0 0 0 io_out[0]
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 8338 0 0 0 io_out[10]
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 8338 0 0 0 io_out[11]
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 8338 0 0 0 io_out[12]
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 8338 0 0 0 io_out[13]
flabel metal3 s -800 506802 480 506914 0 FreeSans 8338 0 0 0 io_out[14]
flabel metal3 s -800 463580 480 463692 0 FreeSans 8338 0 0 0 io_out[15]
flabel metal3 s -800 420358 480 420470 0 FreeSans 8338 0 0 0 io_out[16]
flabel metal3 s -800 377136 480 377248 0 FreeSans 8338 0 0 0 io_out[17]
flabel metal3 s -800 333914 480 334026 0 FreeSans 8338 0 0 0 io_out[18]
flabel metal3 s -800 290692 480 290804 0 FreeSans 8338 0 0 0 io_out[19]
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 8338 0 0 0 io_out[1]
flabel metal3 s -800 247670 480 247782 0 FreeSans 8338 0 0 0 io_out[20]
flabel metal3 s -800 120048 480 120160 0 FreeSans 8338 0 0 0 io_out[21]
flabel metal3 s -800 76826 480 76938 0 FreeSans 8338 0 0 0 io_out[22]
flabel metal3 s -800 33604 480 33716 0 FreeSans 8338 0 0 0 io_out[23]
flabel metal3 s -800 12182 480 12294 0 FreeSans 8338 0 0 0 io_out[24]
flabel metal3 s -800 7454 480 7566 0 FreeSans 8338 0 0 0 io_out[25]
flabel metal3 s -800 2726 480 2838 0 FreeSans 8338 0 0 0 io_out[26]
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 8338 0 0 0 io_out[2]
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 8338 0 0 0 io_out[3]
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 8338 0 0 0 io_out[4]
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 8338 0 0 0 io_out[5]
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 8338 0 0 0 io_out[6]
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 8338 0 0 0 io_out[7]
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 8338 0 0 0 io_out[8]
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 8338 0 0 0 io_out[9]
flabel metal2 s 125816 -800 125928 480 0 FreeSans 8338 90 0 0 la_data_in[0]
flabel metal2 s 480416 -800 480528 480 0 FreeSans 8338 90 0 0 la_data_in[100]
flabel metal2 s 483962 -800 484074 480 0 FreeSans 8338 90 0 0 la_data_in[101]
flabel metal2 s 487508 -800 487620 480 0 FreeSans 8338 90 0 0 la_data_in[102]
flabel metal2 s 491054 -800 491166 480 0 FreeSans 8338 90 0 0 la_data_in[103]
flabel metal2 s 494600 -800 494712 480 0 FreeSans 8338 90 0 0 la_data_in[104]
flabel metal2 s 498146 -800 498258 480 0 FreeSans 8338 90 0 0 la_data_in[105]
flabel metal2 s 501692 -800 501804 480 0 FreeSans 8338 90 0 0 la_data_in[106]
flabel metal2 s 505238 -800 505350 480 0 FreeSans 8338 90 0 0 la_data_in[107]
flabel metal2 s 508784 -800 508896 480 0 FreeSans 8338 90 0 0 la_data_in[108]
flabel metal2 s 512330 -800 512442 480 0 FreeSans 8338 90 0 0 la_data_in[109]
flabel metal2 s 161276 -800 161388 480 0 FreeSans 8338 90 0 0 la_data_in[10]
flabel metal2 s 515876 -800 515988 480 0 FreeSans 8338 90 0 0 la_data_in[110]
flabel metal2 s 519422 -800 519534 480 0 FreeSans 8338 90 0 0 la_data_in[111]
flabel metal2 s 522968 -800 523080 480 0 FreeSans 8338 90 0 0 la_data_in[112]
flabel metal2 s 526514 -800 526626 480 0 FreeSans 8338 90 0 0 la_data_in[113]
flabel metal2 s 530060 -800 530172 480 0 FreeSans 8338 90 0 0 la_data_in[114]
flabel metal2 s 533606 -800 533718 480 0 FreeSans 8338 90 0 0 la_data_in[115]
flabel metal2 s 537152 -800 537264 480 0 FreeSans 8338 90 0 0 la_data_in[116]
flabel metal2 s 540698 -800 540810 480 0 FreeSans 8338 90 0 0 la_data_in[117]
flabel metal2 s 544244 -800 544356 480 0 FreeSans 8338 90 0 0 la_data_in[118]
flabel metal2 s 547790 -800 547902 480 0 FreeSans 8338 90 0 0 la_data_in[119]
flabel metal2 s 164822 -800 164934 480 0 FreeSans 8338 90 0 0 la_data_in[11]
flabel metal2 s 551336 -800 551448 480 0 FreeSans 8338 90 0 0 la_data_in[120]
flabel metal2 s 554882 -800 554994 480 0 FreeSans 8338 90 0 0 la_data_in[121]
flabel metal2 s 558428 -800 558540 480 0 FreeSans 8338 90 0 0 la_data_in[122]
flabel metal2 s 561974 -800 562086 480 0 FreeSans 8338 90 0 0 la_data_in[123]
flabel metal2 s 565520 -800 565632 480 0 FreeSans 8338 90 0 0 la_data_in[124]
flabel metal2 s 569066 -800 569178 480 0 FreeSans 8338 90 0 0 la_data_in[125]
flabel metal2 s 572612 -800 572724 480 0 FreeSans 8338 90 0 0 la_data_in[126]
flabel metal2 s 576158 -800 576270 480 0 FreeSans 8338 90 0 0 la_data_in[127]
flabel metal2 s 168368 -800 168480 480 0 FreeSans 8338 90 0 0 la_data_in[12]
flabel metal2 s 171914 -800 172026 480 0 FreeSans 8338 90 0 0 la_data_in[13]
flabel metal2 s 175460 -800 175572 480 0 FreeSans 8338 90 0 0 la_data_in[14]
flabel metal2 s 179006 -800 179118 480 0 FreeSans 8338 90 0 0 la_data_in[15]
flabel metal2 s 182552 -800 182664 480 0 FreeSans 8338 90 0 0 la_data_in[16]
flabel metal2 s 186098 -800 186210 480 0 FreeSans 8338 90 0 0 la_data_in[17]
flabel metal2 s 189644 -800 189756 480 0 FreeSans 8338 90 0 0 la_data_in[18]
flabel metal2 s 193190 -800 193302 480 0 FreeSans 8338 90 0 0 la_data_in[19]
flabel metal2 s 129362 -800 129474 480 0 FreeSans 8338 90 0 0 la_data_in[1]
flabel metal2 s 196736 -800 196848 480 0 FreeSans 8338 90 0 0 la_data_in[20]
flabel metal2 s 200282 -800 200394 480 0 FreeSans 8338 90 0 0 la_data_in[21]
flabel metal2 s 203828 -800 203940 480 0 FreeSans 8338 90 0 0 la_data_in[22]
flabel metal2 s 207374 -800 207486 480 0 FreeSans 8338 90 0 0 la_data_in[23]
flabel metal2 s 210920 -800 211032 480 0 FreeSans 8338 90 0 0 la_data_in[24]
flabel metal2 s 214466 -800 214578 480 0 FreeSans 8338 90 0 0 la_data_in[25]
flabel metal2 s 218012 -800 218124 480 0 FreeSans 8338 90 0 0 la_data_in[26]
flabel metal2 s 221558 -800 221670 480 0 FreeSans 8338 90 0 0 la_data_in[27]
flabel metal2 s 225104 -800 225216 480 0 FreeSans 8338 90 0 0 la_data_in[28]
flabel metal2 s 228650 -800 228762 480 0 FreeSans 8338 90 0 0 la_data_in[29]
flabel metal2 s 132908 -800 133020 480 0 FreeSans 8338 90 0 0 la_data_in[2]
flabel metal2 s 232196 -800 232308 480 0 FreeSans 8338 90 0 0 la_data_in[30]
flabel metal2 s 235742 -800 235854 480 0 FreeSans 8338 90 0 0 la_data_in[31]
flabel metal2 s 239288 -800 239400 480 0 FreeSans 8338 90 0 0 la_data_in[32]
flabel metal2 s 242834 -800 242946 480 0 FreeSans 8338 90 0 0 la_data_in[33]
flabel metal2 s 246380 -800 246492 480 0 FreeSans 8338 90 0 0 la_data_in[34]
flabel metal2 s 249926 -800 250038 480 0 FreeSans 8338 90 0 0 la_data_in[35]
flabel metal2 s 253472 -800 253584 480 0 FreeSans 8338 90 0 0 la_data_in[36]
flabel metal2 s 257018 -800 257130 480 0 FreeSans 8338 90 0 0 la_data_in[37]
flabel metal2 s 260564 -800 260676 480 0 FreeSans 8338 90 0 0 la_data_in[38]
flabel metal2 s 264110 -800 264222 480 0 FreeSans 8338 90 0 0 la_data_in[39]
flabel metal2 s 136454 -800 136566 480 0 FreeSans 8338 90 0 0 la_data_in[3]
flabel metal2 s 267656 -800 267768 480 0 FreeSans 8338 90 0 0 la_data_in[40]
flabel metal2 s 271202 -800 271314 480 0 FreeSans 8338 90 0 0 la_data_in[41]
flabel metal2 s 274748 -800 274860 480 0 FreeSans 8338 90 0 0 la_data_in[42]
flabel metal2 s 278294 -800 278406 480 0 FreeSans 8338 90 0 0 la_data_in[43]
flabel metal2 s 281840 -800 281952 480 0 FreeSans 8338 90 0 0 la_data_in[44]
flabel metal2 s 285386 -800 285498 480 0 FreeSans 8338 90 0 0 la_data_in[45]
flabel metal2 s 288932 -800 289044 480 0 FreeSans 8338 90 0 0 la_data_in[46]
flabel metal2 s 292478 -800 292590 480 0 FreeSans 8338 90 0 0 la_data_in[47]
flabel metal2 s 296024 -800 296136 480 0 FreeSans 8338 90 0 0 la_data_in[48]
flabel metal2 s 299570 -800 299682 480 0 FreeSans 8338 90 0 0 la_data_in[49]
flabel metal2 s 140000 -800 140112 480 0 FreeSans 8338 90 0 0 la_data_in[4]
flabel metal2 s 303116 -800 303228 480 0 FreeSans 8338 90 0 0 la_data_in[50]
flabel metal2 s 306662 -800 306774 480 0 FreeSans 8338 90 0 0 la_data_in[51]
flabel metal2 s 310208 -800 310320 480 0 FreeSans 8338 90 0 0 la_data_in[52]
flabel metal2 s 313754 -800 313866 480 0 FreeSans 8338 90 0 0 la_data_in[53]
flabel metal2 s 317300 -800 317412 480 0 FreeSans 8338 90 0 0 la_data_in[54]
flabel metal2 s 320846 -800 320958 480 0 FreeSans 8338 90 0 0 la_data_in[55]
flabel metal2 s 324392 -800 324504 480 0 FreeSans 8338 90 0 0 la_data_in[56]
flabel metal2 s 327938 -800 328050 480 0 FreeSans 8338 90 0 0 la_data_in[57]
flabel metal2 s 331484 -800 331596 480 0 FreeSans 8338 90 0 0 la_data_in[58]
flabel metal2 s 335030 -800 335142 480 0 FreeSans 8338 90 0 0 la_data_in[59]
flabel metal2 s 143546 -800 143658 480 0 FreeSans 8338 90 0 0 la_data_in[5]
flabel metal2 s 338576 -800 338688 480 0 FreeSans 8338 90 0 0 la_data_in[60]
flabel metal2 s 342122 -800 342234 480 0 FreeSans 8338 90 0 0 la_data_in[61]
flabel metal2 s 345668 -800 345780 480 0 FreeSans 8338 90 0 0 la_data_in[62]
flabel metal2 s 349214 -800 349326 480 0 FreeSans 8338 90 0 0 la_data_in[63]
flabel metal2 s 352760 -800 352872 480 0 FreeSans 8338 90 0 0 la_data_in[64]
flabel metal2 s 356306 -800 356418 480 0 FreeSans 8338 90 0 0 la_data_in[65]
flabel metal2 s 359852 -800 359964 480 0 FreeSans 8338 90 0 0 la_data_in[66]
flabel metal2 s 363398 -800 363510 480 0 FreeSans 8338 90 0 0 la_data_in[67]
flabel metal2 s 366944 -800 367056 480 0 FreeSans 8338 90 0 0 la_data_in[68]
flabel metal2 s 370490 -800 370602 480 0 FreeSans 8338 90 0 0 la_data_in[69]
flabel metal2 s 147092 -800 147204 480 0 FreeSans 8338 90 0 0 la_data_in[6]
flabel metal2 s 374036 -800 374148 480 0 FreeSans 8338 90 0 0 la_data_in[70]
flabel metal2 s 377582 -800 377694 480 0 FreeSans 8338 90 0 0 la_data_in[71]
flabel metal2 s 381128 -800 381240 480 0 FreeSans 8338 90 0 0 la_data_in[72]
flabel metal2 s 384674 -800 384786 480 0 FreeSans 8338 90 0 0 la_data_in[73]
flabel metal2 s 388220 -800 388332 480 0 FreeSans 8338 90 0 0 la_data_in[74]
flabel metal2 s 391766 -800 391878 480 0 FreeSans 8338 90 0 0 la_data_in[75]
flabel metal2 s 395312 -800 395424 480 0 FreeSans 8338 90 0 0 la_data_in[76]
flabel metal2 s 398858 -800 398970 480 0 FreeSans 8338 90 0 0 la_data_in[77]
flabel metal2 s 402404 -800 402516 480 0 FreeSans 8338 90 0 0 la_data_in[78]
flabel metal2 s 405950 -800 406062 480 0 FreeSans 8338 90 0 0 la_data_in[79]
flabel metal2 s 150638 -800 150750 480 0 FreeSans 8338 90 0 0 la_data_in[7]
flabel metal2 s 409496 -800 409608 480 0 FreeSans 8338 90 0 0 la_data_in[80]
flabel metal2 s 413042 -800 413154 480 0 FreeSans 8338 90 0 0 la_data_in[81]
flabel metal2 s 416588 -800 416700 480 0 FreeSans 8338 90 0 0 la_data_in[82]
flabel metal2 s 420134 -800 420246 480 0 FreeSans 8338 90 0 0 la_data_in[83]
flabel metal2 s 423680 -800 423792 480 0 FreeSans 8338 90 0 0 la_data_in[84]
flabel metal2 s 427226 -800 427338 480 0 FreeSans 8338 90 0 0 la_data_in[85]
flabel metal2 s 430772 -800 430884 480 0 FreeSans 8338 90 0 0 la_data_in[86]
flabel metal2 s 434318 -800 434430 480 0 FreeSans 8338 90 0 0 la_data_in[87]
flabel metal2 s 437864 -800 437976 480 0 FreeSans 8338 90 0 0 la_data_in[88]
flabel metal2 s 441410 -800 441522 480 0 FreeSans 8338 90 0 0 la_data_in[89]
flabel metal2 s 154184 -800 154296 480 0 FreeSans 8338 90 0 0 la_data_in[8]
flabel metal2 s 444956 -800 445068 480 0 FreeSans 8338 90 0 0 la_data_in[90]
flabel metal2 s 448502 -800 448614 480 0 FreeSans 8338 90 0 0 la_data_in[91]
flabel metal2 s 452048 -800 452160 480 0 FreeSans 8338 90 0 0 la_data_in[92]
flabel metal2 s 455594 -800 455706 480 0 FreeSans 8338 90 0 0 la_data_in[93]
flabel metal2 s 459140 -800 459252 480 0 FreeSans 8338 90 0 0 la_data_in[94]
flabel metal2 s 462686 -800 462798 480 0 FreeSans 8338 90 0 0 la_data_in[95]
flabel metal2 s 466232 -800 466344 480 0 FreeSans 8338 90 0 0 la_data_in[96]
flabel metal2 s 469778 -800 469890 480 0 FreeSans 8338 90 0 0 la_data_in[97]
flabel metal2 s 473324 -800 473436 480 0 FreeSans 8338 90 0 0 la_data_in[98]
flabel metal2 s 476870 -800 476982 480 0 FreeSans 8338 90 0 0 la_data_in[99]
flabel metal2 s 157730 -800 157842 480 0 FreeSans 8338 90 0 0 la_data_in[9]
flabel metal2 s 126998 -800 127110 480 0 FreeSans 8338 90 0 0 la_data_out[0]
flabel metal2 s 481598 -800 481710 480 0 FreeSans 8338 90 0 0 la_data_out[100]
flabel metal2 s 485144 -800 485256 480 0 FreeSans 8338 90 0 0 la_data_out[101]
flabel metal2 s 488690 -800 488802 480 0 FreeSans 8338 90 0 0 la_data_out[102]
flabel metal2 s 492236 -800 492348 480 0 FreeSans 8338 90 0 0 la_data_out[103]
flabel metal2 s 495782 -800 495894 480 0 FreeSans 8338 90 0 0 la_data_out[104]
flabel metal2 s 499328 -800 499440 480 0 FreeSans 8338 90 0 0 la_data_out[105]
flabel metal2 s 502874 -800 502986 480 0 FreeSans 8338 90 0 0 la_data_out[106]
flabel metal2 s 506420 -800 506532 480 0 FreeSans 8338 90 0 0 la_data_out[107]
flabel metal2 s 509966 -800 510078 480 0 FreeSans 8338 90 0 0 la_data_out[108]
flabel metal2 s 513512 -800 513624 480 0 FreeSans 8338 90 0 0 la_data_out[109]
flabel metal2 s 162458 -800 162570 480 0 FreeSans 8338 90 0 0 la_data_out[10]
flabel metal2 s 517058 -800 517170 480 0 FreeSans 8338 90 0 0 la_data_out[110]
flabel metal2 s 520604 -800 520716 480 0 FreeSans 8338 90 0 0 la_data_out[111]
flabel metal2 s 524150 -800 524262 480 0 FreeSans 8338 90 0 0 la_data_out[112]
flabel metal2 s 527696 -800 527808 480 0 FreeSans 8338 90 0 0 la_data_out[113]
flabel metal2 s 531242 -800 531354 480 0 FreeSans 8338 90 0 0 la_data_out[114]
flabel metal2 s 534788 -800 534900 480 0 FreeSans 8338 90 0 0 la_data_out[115]
flabel metal2 s 538334 -800 538446 480 0 FreeSans 8338 90 0 0 la_data_out[116]
flabel metal2 s 541880 -800 541992 480 0 FreeSans 8338 90 0 0 la_data_out[117]
flabel metal2 s 545426 -800 545538 480 0 FreeSans 8338 90 0 0 la_data_out[118]
flabel metal2 s 548972 -800 549084 480 0 FreeSans 8338 90 0 0 la_data_out[119]
flabel metal2 s 166004 -800 166116 480 0 FreeSans 8338 90 0 0 la_data_out[11]
flabel metal2 s 552518 -800 552630 480 0 FreeSans 8338 90 0 0 la_data_out[120]
flabel metal2 s 556064 -800 556176 480 0 FreeSans 8338 90 0 0 la_data_out[121]
flabel metal2 s 559610 -800 559722 480 0 FreeSans 8338 90 0 0 la_data_out[122]
flabel metal2 s 563156 -800 563268 480 0 FreeSans 8338 90 0 0 la_data_out[123]
flabel metal2 s 566702 -800 566814 480 0 FreeSans 8338 90 0 0 la_data_out[124]
flabel metal2 s 570248 -800 570360 480 0 FreeSans 8338 90 0 0 la_data_out[125]
flabel metal2 s 573794 -800 573906 480 0 FreeSans 8338 90 0 0 la_data_out[126]
flabel metal2 s 577340 -800 577452 480 0 FreeSans 8338 90 0 0 la_data_out[127]
flabel metal2 s 169550 -800 169662 480 0 FreeSans 8338 90 0 0 la_data_out[12]
flabel metal2 s 173096 -800 173208 480 0 FreeSans 8338 90 0 0 la_data_out[13]
flabel metal2 s 176642 -800 176754 480 0 FreeSans 8338 90 0 0 la_data_out[14]
flabel metal2 s 180188 -800 180300 480 0 FreeSans 8338 90 0 0 la_data_out[15]
flabel metal2 s 183734 -800 183846 480 0 FreeSans 8338 90 0 0 la_data_out[16]
flabel metal2 s 187280 -800 187392 480 0 FreeSans 8338 90 0 0 la_data_out[17]
flabel metal2 s 190826 -800 190938 480 0 FreeSans 8338 90 0 0 la_data_out[18]
flabel metal2 s 194372 -800 194484 480 0 FreeSans 8338 90 0 0 la_data_out[19]
flabel metal2 s 130544 -800 130656 480 0 FreeSans 8338 90 0 0 la_data_out[1]
flabel metal2 s 197918 -800 198030 480 0 FreeSans 8338 90 0 0 la_data_out[20]
flabel metal2 s 201464 -800 201576 480 0 FreeSans 8338 90 0 0 la_data_out[21]
flabel metal2 s 205010 -800 205122 480 0 FreeSans 8338 90 0 0 la_data_out[22]
flabel metal2 s 208556 -800 208668 480 0 FreeSans 8338 90 0 0 la_data_out[23]
flabel metal2 s 212102 -800 212214 480 0 FreeSans 8338 90 0 0 la_data_out[24]
flabel metal2 s 215648 -800 215760 480 0 FreeSans 8338 90 0 0 la_data_out[25]
flabel metal2 s 219194 -800 219306 480 0 FreeSans 8338 90 0 0 la_data_out[26]
flabel metal2 s 222740 -800 222852 480 0 FreeSans 8338 90 0 0 la_data_out[27]
flabel metal2 s 226286 -800 226398 480 0 FreeSans 8338 90 0 0 la_data_out[28]
flabel metal2 s 229832 -800 229944 480 0 FreeSans 8338 90 0 0 la_data_out[29]
flabel metal2 s 134090 -800 134202 480 0 FreeSans 8338 90 0 0 la_data_out[2]
flabel metal2 s 233378 -800 233490 480 0 FreeSans 8338 90 0 0 la_data_out[30]
flabel metal2 s 236924 -800 237036 480 0 FreeSans 8338 90 0 0 la_data_out[31]
flabel metal2 s 240470 -800 240582 480 0 FreeSans 8338 90 0 0 la_data_out[32]
flabel metal2 s 244016 -800 244128 480 0 FreeSans 8338 90 0 0 la_data_out[33]
flabel metal2 s 247562 -800 247674 480 0 FreeSans 8338 90 0 0 la_data_out[34]
flabel metal2 s 251108 -800 251220 480 0 FreeSans 8338 90 0 0 la_data_out[35]
flabel metal2 s 254654 -800 254766 480 0 FreeSans 8338 90 0 0 la_data_out[36]
flabel metal2 s 258200 -800 258312 480 0 FreeSans 8338 90 0 0 la_data_out[37]
flabel metal2 s 261746 -800 261858 480 0 FreeSans 8338 90 0 0 la_data_out[38]
flabel metal2 s 265292 -800 265404 480 0 FreeSans 8338 90 0 0 la_data_out[39]
flabel metal2 s 137636 -800 137748 480 0 FreeSans 8338 90 0 0 la_data_out[3]
flabel metal2 s 268838 -800 268950 480 0 FreeSans 8338 90 0 0 la_data_out[40]
flabel metal2 s 272384 -800 272496 480 0 FreeSans 8338 90 0 0 la_data_out[41]
flabel metal2 s 275930 -800 276042 480 0 FreeSans 8338 90 0 0 la_data_out[42]
flabel metal2 s 279476 -800 279588 480 0 FreeSans 8338 90 0 0 la_data_out[43]
flabel metal2 s 283022 -800 283134 480 0 FreeSans 8338 90 0 0 la_data_out[44]
flabel metal2 s 286568 -800 286680 480 0 FreeSans 8338 90 0 0 la_data_out[45]
flabel metal2 s 290114 -800 290226 480 0 FreeSans 8338 90 0 0 la_data_out[46]
flabel metal2 s 293660 -800 293772 480 0 FreeSans 8338 90 0 0 la_data_out[47]
flabel metal2 s 297206 -800 297318 480 0 FreeSans 8338 90 0 0 la_data_out[48]
flabel metal2 s 300752 -800 300864 480 0 FreeSans 8338 90 0 0 la_data_out[49]
flabel metal2 s 141182 -800 141294 480 0 FreeSans 8338 90 0 0 la_data_out[4]
flabel metal2 s 304298 -800 304410 480 0 FreeSans 8338 90 0 0 la_data_out[50]
flabel metal2 s 307844 -800 307956 480 0 FreeSans 8338 90 0 0 la_data_out[51]
flabel metal2 s 311390 -800 311502 480 0 FreeSans 8338 90 0 0 la_data_out[52]
flabel metal2 s 314936 -800 315048 480 0 FreeSans 8338 90 0 0 la_data_out[53]
flabel metal2 s 318482 -800 318594 480 0 FreeSans 8338 90 0 0 la_data_out[54]
flabel metal2 s 322028 -800 322140 480 0 FreeSans 8338 90 0 0 la_data_out[55]
flabel metal2 s 325574 -800 325686 480 0 FreeSans 8338 90 0 0 la_data_out[56]
flabel metal2 s 329120 -800 329232 480 0 FreeSans 8338 90 0 0 la_data_out[57]
flabel metal2 s 332666 -800 332778 480 0 FreeSans 8338 90 0 0 la_data_out[58]
flabel metal2 s 336212 -800 336324 480 0 FreeSans 8338 90 0 0 la_data_out[59]
flabel metal2 s 144728 -800 144840 480 0 FreeSans 8338 90 0 0 la_data_out[5]
flabel metal2 s 339758 -800 339870 480 0 FreeSans 8338 90 0 0 la_data_out[60]
flabel metal2 s 343304 -800 343416 480 0 FreeSans 8338 90 0 0 la_data_out[61]
flabel metal2 s 346850 -800 346962 480 0 FreeSans 8338 90 0 0 la_data_out[62]
flabel metal2 s 350396 -800 350508 480 0 FreeSans 8338 90 0 0 la_data_out[63]
flabel metal2 s 353942 -800 354054 480 0 FreeSans 8338 90 0 0 la_data_out[64]
flabel metal2 s 357488 -800 357600 480 0 FreeSans 8338 90 0 0 la_data_out[65]
flabel metal2 s 361034 -800 361146 480 0 FreeSans 8338 90 0 0 la_data_out[66]
flabel metal2 s 364580 -800 364692 480 0 FreeSans 8338 90 0 0 la_data_out[67]
flabel metal2 s 368126 -800 368238 480 0 FreeSans 8338 90 0 0 la_data_out[68]
flabel metal2 s 371672 -800 371784 480 0 FreeSans 8338 90 0 0 la_data_out[69]
flabel metal2 s 148274 -800 148386 480 0 FreeSans 8338 90 0 0 la_data_out[6]
flabel metal2 s 375218 -800 375330 480 0 FreeSans 8338 90 0 0 la_data_out[70]
flabel metal2 s 378764 -800 378876 480 0 FreeSans 8338 90 0 0 la_data_out[71]
flabel metal2 s 382310 -800 382422 480 0 FreeSans 8338 90 0 0 la_data_out[72]
flabel metal2 s 385856 -800 385968 480 0 FreeSans 8338 90 0 0 la_data_out[73]
flabel metal2 s 389402 -800 389514 480 0 FreeSans 8338 90 0 0 la_data_out[74]
flabel metal2 s 392948 -800 393060 480 0 FreeSans 8338 90 0 0 la_data_out[75]
flabel metal2 s 396494 -800 396606 480 0 FreeSans 8338 90 0 0 la_data_out[76]
flabel metal2 s 400040 -800 400152 480 0 FreeSans 8338 90 0 0 la_data_out[77]
flabel metal2 s 403586 -800 403698 480 0 FreeSans 8338 90 0 0 la_data_out[78]
flabel metal2 s 407132 -800 407244 480 0 FreeSans 8338 90 0 0 la_data_out[79]
flabel metal2 s 151820 -800 151932 480 0 FreeSans 8338 90 0 0 la_data_out[7]
flabel metal2 s 410678 -800 410790 480 0 FreeSans 8338 90 0 0 la_data_out[80]
flabel metal2 s 414224 -800 414336 480 0 FreeSans 8338 90 0 0 la_data_out[81]
flabel metal2 s 417770 -800 417882 480 0 FreeSans 8338 90 0 0 la_data_out[82]
flabel metal2 s 421316 -800 421428 480 0 FreeSans 8338 90 0 0 la_data_out[83]
flabel metal2 s 424862 -800 424974 480 0 FreeSans 8338 90 0 0 la_data_out[84]
flabel metal2 s 428408 -800 428520 480 0 FreeSans 8338 90 0 0 la_data_out[85]
flabel metal2 s 431954 -800 432066 480 0 FreeSans 8338 90 0 0 la_data_out[86]
flabel metal2 s 435500 -800 435612 480 0 FreeSans 8338 90 0 0 la_data_out[87]
flabel metal2 s 439046 -800 439158 480 0 FreeSans 8338 90 0 0 la_data_out[88]
flabel metal2 s 442592 -800 442704 480 0 FreeSans 8338 90 0 0 la_data_out[89]
flabel metal2 s 155366 -800 155478 480 0 FreeSans 8338 90 0 0 la_data_out[8]
flabel metal2 s 446138 -800 446250 480 0 FreeSans 8338 90 0 0 la_data_out[90]
flabel metal2 s 449684 -800 449796 480 0 FreeSans 8338 90 0 0 la_data_out[91]
flabel metal2 s 453230 -800 453342 480 0 FreeSans 8338 90 0 0 la_data_out[92]
flabel metal2 s 456776 -800 456888 480 0 FreeSans 8338 90 0 0 la_data_out[93]
flabel metal2 s 460322 -800 460434 480 0 FreeSans 8338 90 0 0 la_data_out[94]
flabel metal2 s 463868 -800 463980 480 0 FreeSans 8338 90 0 0 la_data_out[95]
flabel metal2 s 467414 -800 467526 480 0 FreeSans 8338 90 0 0 la_data_out[96]
flabel metal2 s 470960 -800 471072 480 0 FreeSans 8338 90 0 0 la_data_out[97]
flabel metal2 s 474506 -800 474618 480 0 FreeSans 8338 90 0 0 la_data_out[98]
flabel metal2 s 478052 -800 478164 480 0 FreeSans 8338 90 0 0 la_data_out[99]
flabel metal2 s 158912 -800 159024 480 0 FreeSans 8338 90 0 0 la_data_out[9]
flabel metal2 s 128180 -800 128292 480 0 FreeSans 8338 90 0 0 la_oenb[0]
flabel metal2 s 482780 -800 482892 480 0 FreeSans 8338 90 0 0 la_oenb[100]
flabel metal2 s 486326 -800 486438 480 0 FreeSans 8338 90 0 0 la_oenb[101]
flabel metal2 s 489872 -800 489984 480 0 FreeSans 8338 90 0 0 la_oenb[102]
flabel metal2 s 493418 -800 493530 480 0 FreeSans 8338 90 0 0 la_oenb[103]
flabel metal2 s 496964 -800 497076 480 0 FreeSans 8338 90 0 0 la_oenb[104]
flabel metal2 s 500510 -800 500622 480 0 FreeSans 8338 90 0 0 la_oenb[105]
flabel metal2 s 504056 -800 504168 480 0 FreeSans 8338 90 0 0 la_oenb[106]
flabel metal2 s 507602 -800 507714 480 0 FreeSans 8338 90 0 0 la_oenb[107]
flabel metal2 s 511148 -800 511260 480 0 FreeSans 8338 90 0 0 la_oenb[108]
flabel metal2 s 514694 -800 514806 480 0 FreeSans 8338 90 0 0 la_oenb[109]
flabel metal2 s 163640 -800 163752 480 0 FreeSans 8338 90 0 0 la_oenb[10]
flabel metal2 s 518240 -800 518352 480 0 FreeSans 8338 90 0 0 la_oenb[110]
flabel metal2 s 521786 -800 521898 480 0 FreeSans 8338 90 0 0 la_oenb[111]
flabel metal2 s 525332 -800 525444 480 0 FreeSans 8338 90 0 0 la_oenb[112]
flabel metal2 s 528878 -800 528990 480 0 FreeSans 8338 90 0 0 la_oenb[113]
flabel metal2 s 532424 -800 532536 480 0 FreeSans 8338 90 0 0 la_oenb[114]
flabel metal2 s 535970 -800 536082 480 0 FreeSans 8338 90 0 0 la_oenb[115]
flabel metal2 s 539516 -800 539628 480 0 FreeSans 8338 90 0 0 la_oenb[116]
flabel metal2 s 543062 -800 543174 480 0 FreeSans 8338 90 0 0 la_oenb[117]
flabel metal2 s 546608 -800 546720 480 0 FreeSans 8338 90 0 0 la_oenb[118]
flabel metal2 s 550154 -800 550266 480 0 FreeSans 8338 90 0 0 la_oenb[119]
flabel metal2 s 167186 -800 167298 480 0 FreeSans 8338 90 0 0 la_oenb[11]
flabel metal2 s 553700 -800 553812 480 0 FreeSans 8338 90 0 0 la_oenb[120]
flabel metal2 s 557246 -800 557358 480 0 FreeSans 8338 90 0 0 la_oenb[121]
flabel metal2 s 560792 -800 560904 480 0 FreeSans 8338 90 0 0 la_oenb[122]
flabel metal2 s 564338 -800 564450 480 0 FreeSans 8338 90 0 0 la_oenb[123]
flabel metal2 s 567884 -800 567996 480 0 FreeSans 8338 90 0 0 la_oenb[124]
flabel metal2 s 571430 -800 571542 480 0 FreeSans 8338 90 0 0 la_oenb[125]
flabel metal2 s 574976 -800 575088 480 0 FreeSans 8338 90 0 0 la_oenb[126]
flabel metal2 s 578522 -800 578634 480 0 FreeSans 8338 90 0 0 la_oenb[127]
flabel metal2 s 170732 -800 170844 480 0 FreeSans 8338 90 0 0 la_oenb[12]
flabel metal2 s 174278 -800 174390 480 0 FreeSans 8338 90 0 0 la_oenb[13]
flabel metal2 s 177824 -800 177936 480 0 FreeSans 8338 90 0 0 la_oenb[14]
flabel metal2 s 181370 -800 181482 480 0 FreeSans 8338 90 0 0 la_oenb[15]
flabel metal2 s 184916 -800 185028 480 0 FreeSans 8338 90 0 0 la_oenb[16]
flabel metal2 s 188462 -800 188574 480 0 FreeSans 8338 90 0 0 la_oenb[17]
flabel metal2 s 192008 -800 192120 480 0 FreeSans 8338 90 0 0 la_oenb[18]
flabel metal2 s 195554 -800 195666 480 0 FreeSans 8338 90 0 0 la_oenb[19]
flabel metal2 s 131726 -800 131838 480 0 FreeSans 8338 90 0 0 la_oenb[1]
flabel metal2 s 199100 -800 199212 480 0 FreeSans 8338 90 0 0 la_oenb[20]
flabel metal2 s 202646 -800 202758 480 0 FreeSans 8338 90 0 0 la_oenb[21]
flabel metal2 s 206192 -800 206304 480 0 FreeSans 8338 90 0 0 la_oenb[22]
flabel metal2 s 209738 -800 209850 480 0 FreeSans 8338 90 0 0 la_oenb[23]
flabel metal2 s 213284 -800 213396 480 0 FreeSans 8338 90 0 0 la_oenb[24]
flabel metal2 s 216830 -800 216942 480 0 FreeSans 8338 90 0 0 la_oenb[25]
flabel metal2 s 220376 -800 220488 480 0 FreeSans 8338 90 0 0 la_oenb[26]
flabel metal2 s 223922 -800 224034 480 0 FreeSans 8338 90 0 0 la_oenb[27]
flabel metal2 s 227468 -800 227580 480 0 FreeSans 8338 90 0 0 la_oenb[28]
flabel metal2 s 231014 -800 231126 480 0 FreeSans 8338 90 0 0 la_oenb[29]
flabel metal2 s 135272 -800 135384 480 0 FreeSans 8338 90 0 0 la_oenb[2]
flabel metal2 s 234560 -800 234672 480 0 FreeSans 8338 90 0 0 la_oenb[30]
flabel metal2 s 238106 -800 238218 480 0 FreeSans 8338 90 0 0 la_oenb[31]
flabel metal2 s 241652 -800 241764 480 0 FreeSans 8338 90 0 0 la_oenb[32]
flabel metal2 s 245198 -800 245310 480 0 FreeSans 8338 90 0 0 la_oenb[33]
flabel metal2 s 248744 -800 248856 480 0 FreeSans 8338 90 0 0 la_oenb[34]
flabel metal2 s 252290 -800 252402 480 0 FreeSans 8338 90 0 0 la_oenb[35]
flabel metal2 s 255836 -800 255948 480 0 FreeSans 8338 90 0 0 la_oenb[36]
flabel metal2 s 259382 -800 259494 480 0 FreeSans 8338 90 0 0 la_oenb[37]
flabel metal2 s 262928 -800 263040 480 0 FreeSans 8338 90 0 0 la_oenb[38]
flabel metal2 s 266474 -800 266586 480 0 FreeSans 8338 90 0 0 la_oenb[39]
flabel metal2 s 138818 -800 138930 480 0 FreeSans 8338 90 0 0 la_oenb[3]
flabel metal2 s 270020 -800 270132 480 0 FreeSans 8338 90 0 0 la_oenb[40]
flabel metal2 s 273566 -800 273678 480 0 FreeSans 8338 90 0 0 la_oenb[41]
flabel metal2 s 277112 -800 277224 480 0 FreeSans 8338 90 0 0 la_oenb[42]
flabel metal2 s 280658 -800 280770 480 0 FreeSans 8338 90 0 0 la_oenb[43]
flabel metal2 s 284204 -800 284316 480 0 FreeSans 8338 90 0 0 la_oenb[44]
flabel metal2 s 287750 -800 287862 480 0 FreeSans 8338 90 0 0 la_oenb[45]
flabel metal2 s 291296 -800 291408 480 0 FreeSans 8338 90 0 0 la_oenb[46]
flabel metal2 s 294842 -800 294954 480 0 FreeSans 8338 90 0 0 la_oenb[47]
flabel metal2 s 298388 -800 298500 480 0 FreeSans 8338 90 0 0 la_oenb[48]
flabel metal2 s 301934 -800 302046 480 0 FreeSans 8338 90 0 0 la_oenb[49]
flabel metal2 s 142364 -800 142476 480 0 FreeSans 8338 90 0 0 la_oenb[4]
flabel metal2 s 305480 -800 305592 480 0 FreeSans 8338 90 0 0 la_oenb[50]
flabel metal2 s 309026 -800 309138 480 0 FreeSans 8338 90 0 0 la_oenb[51]
flabel metal2 s 312572 -800 312684 480 0 FreeSans 8338 90 0 0 la_oenb[52]
flabel metal2 s 316118 -800 316230 480 0 FreeSans 8338 90 0 0 la_oenb[53]
flabel metal2 s 319664 -800 319776 480 0 FreeSans 8338 90 0 0 la_oenb[54]
flabel metal2 s 323210 -800 323322 480 0 FreeSans 8338 90 0 0 la_oenb[55]
flabel metal2 s 326756 -800 326868 480 0 FreeSans 8338 90 0 0 la_oenb[56]
flabel metal2 s 330302 -800 330414 480 0 FreeSans 8338 90 0 0 la_oenb[57]
flabel metal2 s 333848 -800 333960 480 0 FreeSans 8338 90 0 0 la_oenb[58]
flabel metal2 s 337394 -800 337506 480 0 FreeSans 8338 90 0 0 la_oenb[59]
flabel metal2 s 145910 -800 146022 480 0 FreeSans 8338 90 0 0 la_oenb[5]
flabel metal2 s 340940 -800 341052 480 0 FreeSans 8338 90 0 0 la_oenb[60]
flabel metal2 s 344486 -800 344598 480 0 FreeSans 8338 90 0 0 la_oenb[61]
flabel metal2 s 348032 -800 348144 480 0 FreeSans 8338 90 0 0 la_oenb[62]
flabel metal2 s 351578 -800 351690 480 0 FreeSans 8338 90 0 0 la_oenb[63]
flabel metal2 s 355124 -800 355236 480 0 FreeSans 8338 90 0 0 la_oenb[64]
flabel metal2 s 358670 -800 358782 480 0 FreeSans 8338 90 0 0 la_oenb[65]
flabel metal2 s 362216 -800 362328 480 0 FreeSans 8338 90 0 0 la_oenb[66]
flabel metal2 s 365762 -800 365874 480 0 FreeSans 8338 90 0 0 la_oenb[67]
flabel metal2 s 369308 -800 369420 480 0 FreeSans 8338 90 0 0 la_oenb[68]
flabel metal2 s 372854 -800 372966 480 0 FreeSans 8338 90 0 0 la_oenb[69]
flabel metal2 s 149456 -800 149568 480 0 FreeSans 8338 90 0 0 la_oenb[6]
flabel metal2 s 376400 -800 376512 480 0 FreeSans 8338 90 0 0 la_oenb[70]
flabel metal2 s 379946 -800 380058 480 0 FreeSans 8338 90 0 0 la_oenb[71]
flabel metal2 s 383492 -800 383604 480 0 FreeSans 8338 90 0 0 la_oenb[72]
flabel metal2 s 387038 -800 387150 480 0 FreeSans 8338 90 0 0 la_oenb[73]
flabel metal2 s 390584 -800 390696 480 0 FreeSans 8338 90 0 0 la_oenb[74]
flabel metal2 s 394130 -800 394242 480 0 FreeSans 8338 90 0 0 la_oenb[75]
flabel metal2 s 397676 -800 397788 480 0 FreeSans 8338 90 0 0 la_oenb[76]
flabel metal2 s 401222 -800 401334 480 0 FreeSans 8338 90 0 0 la_oenb[77]
flabel metal2 s 404768 -800 404880 480 0 FreeSans 8338 90 0 0 la_oenb[78]
flabel metal2 s 408314 -800 408426 480 0 FreeSans 8338 90 0 0 la_oenb[79]
flabel metal2 s 153002 -800 153114 480 0 FreeSans 8338 90 0 0 la_oenb[7]
flabel metal2 s 411860 -800 411972 480 0 FreeSans 8338 90 0 0 la_oenb[80]
flabel metal2 s 415406 -800 415518 480 0 FreeSans 8338 90 0 0 la_oenb[81]
flabel metal2 s 418952 -800 419064 480 0 FreeSans 8338 90 0 0 la_oenb[82]
flabel metal2 s 422498 -800 422610 480 0 FreeSans 8338 90 0 0 la_oenb[83]
flabel metal2 s 426044 -800 426156 480 0 FreeSans 8338 90 0 0 la_oenb[84]
flabel metal2 s 429590 -800 429702 480 0 FreeSans 8338 90 0 0 la_oenb[85]
flabel metal2 s 433136 -800 433248 480 0 FreeSans 8338 90 0 0 la_oenb[86]
flabel metal2 s 436682 -800 436794 480 0 FreeSans 8338 90 0 0 la_oenb[87]
flabel metal2 s 440228 -800 440340 480 0 FreeSans 8338 90 0 0 la_oenb[88]
flabel metal2 s 443774 -800 443886 480 0 FreeSans 8338 90 0 0 la_oenb[89]
flabel metal2 s 156548 -800 156660 480 0 FreeSans 8338 90 0 0 la_oenb[8]
flabel metal2 s 447320 -800 447432 480 0 FreeSans 8338 90 0 0 la_oenb[90]
flabel metal2 s 450866 -800 450978 480 0 FreeSans 8338 90 0 0 la_oenb[91]
flabel metal2 s 454412 -800 454524 480 0 FreeSans 8338 90 0 0 la_oenb[92]
flabel metal2 s 457958 -800 458070 480 0 FreeSans 8338 90 0 0 la_oenb[93]
flabel metal2 s 461504 -800 461616 480 0 FreeSans 8338 90 0 0 la_oenb[94]
flabel metal2 s 465050 -800 465162 480 0 FreeSans 8338 90 0 0 la_oenb[95]
flabel metal2 s 468596 -800 468708 480 0 FreeSans 8338 90 0 0 la_oenb[96]
flabel metal2 s 472142 -800 472254 480 0 FreeSans 8338 90 0 0 la_oenb[97]
flabel metal2 s 475688 -800 475800 480 0 FreeSans 8338 90 0 0 la_oenb[98]
flabel metal2 s 479234 -800 479346 480 0 FreeSans 8338 90 0 0 la_oenb[99]
flabel metal2 s 160094 -800 160206 480 0 FreeSans 8338 90 0 0 la_oenb[9]
flabel metal2 s 579704 -800 579816 480 0 FreeSans 8338 90 0 0 user_clock2
flabel metal2 s 580886 -800 580998 480 0 FreeSans 8338 90 0 0 user_irq[0]
flabel metal2 s 582068 -800 582180 480 0 FreeSans 8338 90 0 0 user_irq[1]
flabel metal2 s 583250 -800 583362 480 0 FreeSans 8338 90 0 0 user_irq[2]
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 8338 0 0 0 vccd1
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 8338 0 0 0 vccd1
flabel metal3 s 0 643842 1660 648642 0 FreeSans 8338 0 0 0 vccd2
flabel metal3 s 0 633842 1660 638642 0 FreeSans 8338 0 0 0 vccd2
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 8338 0 0 0 vdda1
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 8338 0 0 0 vdda1
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 8338 0 0 0 vdda1
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 8338 0 0 0 vdda1
flabel metal3 s 0 204888 1660 209688 0 FreeSans 8338 0 0 0 vdda2
flabel metal3 s 0 214888 1660 219688 0 FreeSans 8338 0 0 0 vdda2
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 14300 180 0 0 vssa1
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 14300 180 0 0 vssa1
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 8338 0 0 0 vssa1
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 8338 0 0 0 vssa1
flabel metal3 s 0 559442 1660 564242 0 FreeSans 8338 0 0 0 vssa2
flabel metal3 s 0 549442 1660 554242 0 FreeSans 8338 0 0 0 vssa2
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 8338 0 0 0 vssd1
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 8338 0 0 0 vssd1
flabel metal3 s 0 172888 1660 177688 0 FreeSans 8338 0 0 0 vssd2
flabel metal3 s 0 162888 1660 167688 0 FreeSans 8338 0 0 0 vssd2
flabel metal2 s 524 -800 636 480 0 FreeSans 8338 90 0 0 wb_clk_i
flabel metal2 s 1706 -800 1818 480 0 FreeSans 8338 90 0 0 wb_rst_i
flabel metal2 s 2888 -800 3000 480 0 FreeSans 8338 90 0 0 wbs_ack_o
flabel metal2 s 7616 -800 7728 480 0 FreeSans 8338 90 0 0 wbs_adr_i[0]
flabel metal2 s 47804 -800 47916 480 0 FreeSans 8338 90 0 0 wbs_adr_i[10]
flabel metal2 s 51350 -800 51462 480 0 FreeSans 8338 90 0 0 wbs_adr_i[11]
flabel metal2 s 54896 -800 55008 480 0 FreeSans 8338 90 0 0 wbs_adr_i[12]
flabel metal2 s 58442 -800 58554 480 0 FreeSans 8338 90 0 0 wbs_adr_i[13]
flabel metal2 s 61988 -800 62100 480 0 FreeSans 8338 90 0 0 wbs_adr_i[14]
flabel metal2 s 65534 -800 65646 480 0 FreeSans 8338 90 0 0 wbs_adr_i[15]
flabel metal2 s 69080 -800 69192 480 0 FreeSans 8338 90 0 0 wbs_adr_i[16]
flabel metal2 s 72626 -800 72738 480 0 FreeSans 8338 90 0 0 wbs_adr_i[17]
flabel metal2 s 76172 -800 76284 480 0 FreeSans 8338 90 0 0 wbs_adr_i[18]
flabel metal2 s 79718 -800 79830 480 0 FreeSans 8338 90 0 0 wbs_adr_i[19]
flabel metal2 s 12344 -800 12456 480 0 FreeSans 8338 90 0 0 wbs_adr_i[1]
flabel metal2 s 83264 -800 83376 480 0 FreeSans 8338 90 0 0 wbs_adr_i[20]
flabel metal2 s 86810 -800 86922 480 0 FreeSans 8338 90 0 0 wbs_adr_i[21]
flabel metal2 s 90356 -800 90468 480 0 FreeSans 8338 90 0 0 wbs_adr_i[22]
flabel metal2 s 93902 -800 94014 480 0 FreeSans 8338 90 0 0 wbs_adr_i[23]
flabel metal2 s 97448 -800 97560 480 0 FreeSans 8338 90 0 0 wbs_adr_i[24]
flabel metal2 s 100994 -800 101106 480 0 FreeSans 8338 90 0 0 wbs_adr_i[25]
flabel metal2 s 104540 -800 104652 480 0 FreeSans 8338 90 0 0 wbs_adr_i[26]
flabel metal2 s 108086 -800 108198 480 0 FreeSans 8338 90 0 0 wbs_adr_i[27]
flabel metal2 s 111632 -800 111744 480 0 FreeSans 8338 90 0 0 wbs_adr_i[28]
flabel metal2 s 115178 -800 115290 480 0 FreeSans 8338 90 0 0 wbs_adr_i[29]
flabel metal2 s 17072 -800 17184 480 0 FreeSans 8338 90 0 0 wbs_adr_i[2]
flabel metal2 s 118724 -800 118836 480 0 FreeSans 8338 90 0 0 wbs_adr_i[30]
flabel metal2 s 122270 -800 122382 480 0 FreeSans 8338 90 0 0 wbs_adr_i[31]
flabel metal2 s 21800 -800 21912 480 0 FreeSans 8338 90 0 0 wbs_adr_i[3]
flabel metal2 s 26528 -800 26640 480 0 FreeSans 8338 90 0 0 wbs_adr_i[4]
flabel metal2 s 30074 -800 30186 480 0 FreeSans 8338 90 0 0 wbs_adr_i[5]
flabel metal2 s 33620 -800 33732 480 0 FreeSans 8338 90 0 0 wbs_adr_i[6]
flabel metal2 s 37166 -800 37278 480 0 FreeSans 8338 90 0 0 wbs_adr_i[7]
flabel metal2 s 40712 -800 40824 480 0 FreeSans 8338 90 0 0 wbs_adr_i[8]
flabel metal2 s 44258 -800 44370 480 0 FreeSans 8338 90 0 0 wbs_adr_i[9]
flabel metal2 s 4070 -800 4182 480 0 FreeSans 8338 90 0 0 wbs_cyc_i
flabel metal2 s 8798 -800 8910 480 0 FreeSans 8338 90 0 0 wbs_dat_i[0]
flabel metal2 s 48986 -800 49098 480 0 FreeSans 8338 90 0 0 wbs_dat_i[10]
flabel metal2 s 52532 -800 52644 480 0 FreeSans 8338 90 0 0 wbs_dat_i[11]
flabel metal2 s 56078 -800 56190 480 0 FreeSans 8338 90 0 0 wbs_dat_i[12]
flabel metal2 s 59624 -800 59736 480 0 FreeSans 8338 90 0 0 wbs_dat_i[13]
flabel metal2 s 63170 -800 63282 480 0 FreeSans 8338 90 0 0 wbs_dat_i[14]
flabel metal2 s 66716 -800 66828 480 0 FreeSans 8338 90 0 0 wbs_dat_i[15]
flabel metal2 s 70262 -800 70374 480 0 FreeSans 8338 90 0 0 wbs_dat_i[16]
flabel metal2 s 73808 -800 73920 480 0 FreeSans 8338 90 0 0 wbs_dat_i[17]
flabel metal2 s 77354 -800 77466 480 0 FreeSans 8338 90 0 0 wbs_dat_i[18]
flabel metal2 s 80900 -800 81012 480 0 FreeSans 8338 90 0 0 wbs_dat_i[19]
flabel metal2 s 13526 -800 13638 480 0 FreeSans 8338 90 0 0 wbs_dat_i[1]
flabel metal2 s 84446 -800 84558 480 0 FreeSans 8338 90 0 0 wbs_dat_i[20]
flabel metal2 s 87992 -800 88104 480 0 FreeSans 8338 90 0 0 wbs_dat_i[21]
flabel metal2 s 91538 -800 91650 480 0 FreeSans 8338 90 0 0 wbs_dat_i[22]
flabel metal2 s 95084 -800 95196 480 0 FreeSans 8338 90 0 0 wbs_dat_i[23]
flabel metal2 s 98630 -800 98742 480 0 FreeSans 8338 90 0 0 wbs_dat_i[24]
flabel metal2 s 102176 -800 102288 480 0 FreeSans 8338 90 0 0 wbs_dat_i[25]
flabel metal2 s 105722 -800 105834 480 0 FreeSans 8338 90 0 0 wbs_dat_i[26]
flabel metal2 s 109268 -800 109380 480 0 FreeSans 8338 90 0 0 wbs_dat_i[27]
flabel metal2 s 112814 -800 112926 480 0 FreeSans 8338 90 0 0 wbs_dat_i[28]
flabel metal2 s 116360 -800 116472 480 0 FreeSans 8338 90 0 0 wbs_dat_i[29]
flabel metal2 s 18254 -800 18366 480 0 FreeSans 8338 90 0 0 wbs_dat_i[2]
flabel metal2 s 119906 -800 120018 480 0 FreeSans 8338 90 0 0 wbs_dat_i[30]
flabel metal2 s 123452 -800 123564 480 0 FreeSans 8338 90 0 0 wbs_dat_i[31]
flabel metal2 s 22982 -800 23094 480 0 FreeSans 8338 90 0 0 wbs_dat_i[3]
flabel metal2 s 27710 -800 27822 480 0 FreeSans 8338 90 0 0 wbs_dat_i[4]
flabel metal2 s 31256 -800 31368 480 0 FreeSans 8338 90 0 0 wbs_dat_i[5]
flabel metal2 s 34802 -800 34914 480 0 FreeSans 8338 90 0 0 wbs_dat_i[6]
flabel metal2 s 38348 -800 38460 480 0 FreeSans 8338 90 0 0 wbs_dat_i[7]
flabel metal2 s 41894 -800 42006 480 0 FreeSans 8338 90 0 0 wbs_dat_i[8]
flabel metal2 s 45440 -800 45552 480 0 FreeSans 8338 90 0 0 wbs_dat_i[9]
flabel metal2 s 9980 -800 10092 480 0 FreeSans 8338 90 0 0 wbs_dat_o[0]
flabel metal2 s 50168 -800 50280 480 0 FreeSans 8338 90 0 0 wbs_dat_o[10]
flabel metal2 s 53714 -800 53826 480 0 FreeSans 8338 90 0 0 wbs_dat_o[11]
flabel metal2 s 57260 -800 57372 480 0 FreeSans 8338 90 0 0 wbs_dat_o[12]
flabel metal2 s 60806 -800 60918 480 0 FreeSans 8338 90 0 0 wbs_dat_o[13]
flabel metal2 s 64352 -800 64464 480 0 FreeSans 8338 90 0 0 wbs_dat_o[14]
flabel metal2 s 67898 -800 68010 480 0 FreeSans 8338 90 0 0 wbs_dat_o[15]
flabel metal2 s 71444 -800 71556 480 0 FreeSans 8338 90 0 0 wbs_dat_o[16]
flabel metal2 s 74990 -800 75102 480 0 FreeSans 8338 90 0 0 wbs_dat_o[17]
flabel metal2 s 78536 -800 78648 480 0 FreeSans 8338 90 0 0 wbs_dat_o[18]
flabel metal2 s 82082 -800 82194 480 0 FreeSans 8338 90 0 0 wbs_dat_o[19]
flabel metal2 s 14708 -800 14820 480 0 FreeSans 8338 90 0 0 wbs_dat_o[1]
flabel metal2 s 85628 -800 85740 480 0 FreeSans 8338 90 0 0 wbs_dat_o[20]
flabel metal2 s 89174 -800 89286 480 0 FreeSans 8338 90 0 0 wbs_dat_o[21]
flabel metal2 s 92720 -800 92832 480 0 FreeSans 8338 90 0 0 wbs_dat_o[22]
flabel metal2 s 96266 -800 96378 480 0 FreeSans 8338 90 0 0 wbs_dat_o[23]
flabel metal2 s 99812 -800 99924 480 0 FreeSans 8338 90 0 0 wbs_dat_o[24]
flabel metal2 s 103358 -800 103470 480 0 FreeSans 8338 90 0 0 wbs_dat_o[25]
flabel metal2 s 106904 -800 107016 480 0 FreeSans 8338 90 0 0 wbs_dat_o[26]
flabel metal2 s 110450 -800 110562 480 0 FreeSans 8338 90 0 0 wbs_dat_o[27]
flabel metal2 s 113996 -800 114108 480 0 FreeSans 8338 90 0 0 wbs_dat_o[28]
flabel metal2 s 117542 -800 117654 480 0 FreeSans 8338 90 0 0 wbs_dat_o[29]
flabel metal2 s 19436 -800 19548 480 0 FreeSans 8338 90 0 0 wbs_dat_o[2]
flabel metal2 s 121088 -800 121200 480 0 FreeSans 8338 90 0 0 wbs_dat_o[30]
flabel metal2 s 124634 -800 124746 480 0 FreeSans 8338 90 0 0 wbs_dat_o[31]
flabel metal2 s 24164 -800 24276 480 0 FreeSans 8338 90 0 0 wbs_dat_o[3]
flabel metal2 s 28892 -800 29004 480 0 FreeSans 8338 90 0 0 wbs_dat_o[4]
flabel metal2 s 32438 -800 32550 480 0 FreeSans 8338 90 0 0 wbs_dat_o[5]
flabel metal2 s 35984 -800 36096 480 0 FreeSans 8338 90 0 0 wbs_dat_o[6]
flabel metal2 s 39530 -800 39642 480 0 FreeSans 8338 90 0 0 wbs_dat_o[7]
flabel metal2 s 43076 -800 43188 480 0 FreeSans 8338 90 0 0 wbs_dat_o[8]
flabel metal2 s 46622 -800 46734 480 0 FreeSans 8338 90 0 0 wbs_dat_o[9]
flabel metal2 s 11162 -800 11274 480 0 FreeSans 8338 90 0 0 wbs_sel_i[0]
flabel metal2 s 15890 -800 16002 480 0 FreeSans 8338 90 0 0 wbs_sel_i[1]
flabel metal2 s 20618 -800 20730 480 0 FreeSans 8338 90 0 0 wbs_sel_i[2]
flabel metal2 s 25346 -800 25458 480 0 FreeSans 8338 90 0 0 wbs_sel_i[3]
flabel metal2 s 5252 -800 5364 480 0 FreeSans 8338 90 0 0 wbs_stb_i
flabel metal2 s 6434 -800 6546 480 0 FreeSans 8338 90 0 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
