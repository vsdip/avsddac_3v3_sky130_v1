magic
tech sky130A
timestamp 1616566027
<< locali >>
rect 398 26957 426 27017
rect 99350 14678 102371 14709
rect 97829 14590 98071 14627
rect 97829 14454 97871 14590
rect 97829 14431 97841 14454
rect 97861 14431 97871 14454
rect 97829 14424 97871 14431
rect 97832 14307 97867 14319
rect 97832 14284 97840 14307
rect 97860 14284 97867 14307
rect 97832 11009 97867 14284
rect 102337 12439 102371 14678
rect 102336 12401 102371 12439
rect 97832 10983 97872 11009
rect 82986 2580 83014 2639
rect 83075 2401 83118 2486
rect 83075 2384 83089 2401
rect 83108 2384 83118 2401
rect 83075 2383 83118 2384
rect 84889 1000 84906 1018
rect 84889 995 84913 1000
rect 83074 975 83121 981
rect 83074 964 83087 975
rect 83073 958 83087 964
rect 83106 958 83121 975
rect 83073 948 83121 958
rect 83073 606 83115 948
rect 83069 600 83115 606
rect 84889 603 84906 995
rect 86569 639 86614 1117
rect 86569 612 86577 639
rect 86600 612 86614 639
rect 83069 582 83075 600
rect 83092 582 83115 600
rect 83069 581 83115 582
rect 83070 580 83115 581
rect 84887 597 84916 603
rect 86569 601 86614 612
rect 88277 623 88306 1199
rect 89695 1038 89725 1301
rect 89695 994 89733 1038
rect 88277 601 88284 623
rect 88302 601 88306 623
rect 84887 580 84893 597
rect 84910 580 84916 597
rect 88277 596 88306 601
rect 89697 615 89733 994
rect 89697 592 89707 615
rect 89728 592 89733 615
rect 89697 585 89733 592
rect 91369 617 91394 1383
rect 91369 598 91374 617
rect 91391 598 91394 617
rect 91369 590 91394 598
rect 93988 623 94023 1481
rect 93988 598 93996 623
rect 94018 598 94023 623
rect 93988 588 94023 598
rect 83070 579 83104 580
rect 84887 575 84916 580
rect 83394 507 83430 511
rect 84885 509 84914 516
rect 95734 514 95768 562
rect 83277 501 83435 507
rect 83069 470 83073 489
rect 83090 470 83093 489
rect 83277 478 83402 501
rect 83424 478 83435 501
rect 84885 492 84890 509
rect 84908 492 84914 509
rect 84885 486 84914 492
rect 89701 507 89737 514
rect 83277 471 83435 478
rect 83069 462 83093 470
rect 83069 134 83090 462
rect 83279 285 83299 471
rect 83394 470 83430 471
rect 84888 453 84906 486
rect 89701 484 89709 507
rect 89730 484 89737 507
rect 93986 500 94021 511
rect 88277 473 88310 484
rect 84808 433 84906 453
rect 84810 379 84838 433
rect 84888 431 84906 433
rect 86566 444 86608 466
rect 86566 417 86575 444
rect 86598 417 86608 444
rect 84810 356 84839 379
rect 83279 265 83301 285
rect 83061 111 83090 134
rect 184 -1339 58260 -1335
rect 83061 -1339 83085 111
rect 83281 -959 83301 265
rect 84812 3 84839 356
rect 84812 -17 84840 3
rect 84813 -373 84840 -17
rect 84813 -393 84841 -373
rect 84814 -728 84841 -393
rect 86566 -458 86608 417
rect 84813 -769 84841 -728
rect 86565 -503 86608 -458
rect 88277 451 88284 473
rect 88302 451 88310 473
rect 83281 -973 83305 -959
rect 184 -1358 83085 -1339
rect 184 -1360 58260 -1358
rect 184 -1886 212 -1360
rect 83284 -1409 83305 -973
rect 83279 -1420 83315 -1409
rect 83279 -1445 83284 -1420
rect 83306 -1445 83315 -1420
rect 83279 -1450 83315 -1445
rect 84813 -1433 84840 -769
rect 86565 -1384 86604 -503
rect 86565 -1411 86575 -1384
rect 86598 -1411 86604 -1384
rect 86565 -1420 86604 -1411
rect 88277 -1385 88310 451
rect 89701 104 89737 484
rect 89699 61 89737 104
rect 91370 475 91394 486
rect 91370 456 91374 475
rect 91391 456 91394 475
rect 89699 -405 89731 61
rect 88277 -1412 88281 -1385
rect 88305 -1412 88310 -1385
rect 88277 -1421 88310 -1412
rect 89697 -443 89731 -405
rect 89697 -1372 89729 -443
rect 89697 -1395 89704 -1372
rect 89725 -1395 89729 -1372
rect 89697 -1418 89729 -1395
rect 91370 -1406 91394 456
rect 91369 -1407 91394 -1406
rect 91369 -1426 91373 -1407
rect 91390 -1426 91394 -1407
rect 91369 -1432 91394 -1426
rect 84813 -1454 84816 -1433
rect 84838 -1454 84840 -1433
rect 91370 -1440 91394 -1432
rect 93986 475 93994 500
rect 94016 475 94021 500
rect 93986 -1421 94021 475
rect 93986 -1446 93993 -1421
rect 94015 -1446 94021 -1421
rect 95731 -1403 95768 514
rect 95731 -1429 95736 -1403
rect 95760 -1429 95768 -1403
rect 95731 -1437 95768 -1429
rect 97834 -1428 97872 10983
rect 102336 95 102370 12401
rect 102431 -47 102528 -37
rect 102431 -66 102435 -47
rect 102454 -66 102528 -47
rect 102431 -72 102528 -66
rect 101181 -154 101292 -106
rect 102349 -498 102383 -276
rect 93986 -1454 94021 -1446
rect 97834 -1451 97843 -1428
rect 97864 -1451 97872 -1428
rect 84813 -1458 84840 -1454
rect 97834 -1463 97872 -1451
rect 102027 -527 102383 -498
rect 102027 -530 102377 -527
rect 97831 -1549 97869 -1539
rect 97831 -1572 97841 -1549
rect 97862 -1572 97869 -1549
rect 95724 -1607 95759 -1601
rect 95724 -1633 95730 -1607
rect 95754 -1633 95759 -1607
rect 93985 -1800 94019 -1795
rect 84808 -1824 84846 -1816
rect 84808 -1845 84814 -1824
rect 84836 -1845 84846 -1824
rect 84808 -1851 84846 -1845
rect 86564 -1840 86604 -1813
rect 91372 -1824 91395 -1807
rect 83280 -2227 83303 -2226
rect 83275 -2230 83309 -2227
rect 83275 -2245 83283 -2230
rect 83276 -2247 83283 -2245
rect 83301 -2247 83309 -2230
rect 83276 -2253 83309 -2247
rect 83283 -2501 83300 -2253
rect 84810 -2368 84837 -1851
rect 86564 -1867 86576 -1840
rect 86599 -1867 86604 -1840
rect 84809 -2375 84839 -2368
rect 84809 -2394 84817 -2375
rect 84835 -2394 84839 -2375
rect 84809 -2397 84839 -2394
rect 84812 -2472 84842 -2471
rect 84811 -2476 84842 -2472
rect 84811 -2496 84816 -2476
rect 84837 -2496 84842 -2476
rect 83283 -2510 83301 -2501
rect 84811 -2503 84842 -2496
rect 83283 -2511 83302 -2510
rect 83283 -2518 83300 -2511
rect 84812 -2768 84839 -2503
rect 86564 -2642 86604 -1867
rect 88274 -1840 88307 -1833
rect 88274 -1867 88280 -1840
rect 88304 -1867 88307 -1840
rect 86567 -3307 86601 -2762
rect 88274 -3142 88307 -1867
rect 89699 -1853 89731 -1829
rect 89699 -1876 89704 -1853
rect 89725 -1876 89731 -1853
rect 89699 -2231 89731 -1876
rect 91372 -1843 91374 -1824
rect 91391 -1843 91395 -1824
rect 89699 -2376 89733 -2231
rect 89701 -2754 89733 -2376
rect 89701 -2778 89735 -2754
rect 88274 -3169 88278 -3142
rect 88302 -3169 88307 -3142
rect 88274 -3178 88307 -3169
rect 89703 -3268 89735 -2778
rect 89701 -3301 89735 -3268
rect 86567 -3308 86624 -3307
rect 86567 -3328 86601 -3308
rect 88277 -3377 88313 -3366
rect 88277 -3403 88283 -3377
rect 88306 -3403 88313 -3377
rect 88277 -4938 88313 -3403
rect 89701 -4803 89733 -3301
rect 91372 -3479 91395 -1843
rect 93985 -1825 93993 -1800
rect 94015 -1825 94019 -1800
rect 91372 -3505 91401 -3479
rect 89701 -4826 89707 -4803
rect 89728 -4826 89733 -4803
rect 89701 -4830 89733 -4826
rect 89700 -4919 89735 -4915
rect 89700 -4942 89708 -4919
rect 89729 -4942 89735 -4919
rect 89700 -4948 89735 -4942
rect 89701 -4978 89735 -4948
rect 89703 -5976 89735 -4978
rect 89701 -6002 89735 -5976
rect 89701 -7554 89733 -6002
rect 91374 -7402 91401 -3505
rect 91374 -7409 91405 -7402
rect 91374 -7426 91381 -7409
rect 91398 -7426 91405 -7409
rect 91374 -7431 91405 -7426
rect 91374 -7525 91399 -7524
rect 91371 -7531 91401 -7525
rect 91371 -7548 91376 -7531
rect 91393 -7548 91401 -7531
rect 91371 -7554 91401 -7548
rect 91374 -7911 91399 -7554
rect 91374 -11858 91401 -7911
rect 91374 -11887 91403 -11858
rect 91376 -13860 91403 -11887
rect 93985 -13215 94019 -1825
rect 93985 -13632 94024 -13215
rect 95724 -13863 95759 -1633
rect 97831 -14011 97869 -1572
rect 97832 -14202 97869 -14011
rect 102027 -14137 102054 -530
rect 99148 -14168 102054 -14137
rect 102027 -14169 102054 -14168
rect 97832 -14203 97889 -14202
rect 97832 -14244 97869 -14203
rect 82780 -26291 82810 -26219
<< viali >>
rect 97841 14431 97861 14454
rect 97840 14284 97860 14307
rect 83089 2384 83108 2401
rect 83087 958 83106 975
rect 86577 612 86600 639
rect 83075 582 83092 600
rect 88284 601 88302 623
rect 84893 580 84910 597
rect 89707 592 89728 615
rect 91374 598 91391 617
rect 93996 598 94018 623
rect 83073 470 83090 489
rect 83402 478 83424 501
rect 84890 492 84908 509
rect 89709 484 89730 507
rect 86575 417 86598 444
rect 88284 451 88302 473
rect 83284 -1445 83306 -1420
rect 86575 -1411 86598 -1384
rect 91374 456 91391 475
rect 88281 -1412 88305 -1385
rect 89704 -1395 89725 -1372
rect 91373 -1426 91390 -1407
rect 84816 -1454 84838 -1433
rect 93994 475 94016 500
rect 93993 -1446 94015 -1421
rect 95736 -1429 95760 -1403
rect 102435 -66 102454 -47
rect 97843 -1451 97864 -1428
rect 97841 -1572 97862 -1549
rect 95730 -1633 95754 -1607
rect 84814 -1845 84836 -1824
rect 83283 -2247 83301 -2230
rect 86576 -1867 86599 -1840
rect 84817 -2394 84835 -2375
rect 84816 -2496 84837 -2476
rect 88280 -1867 88304 -1840
rect 89704 -1876 89725 -1853
rect 91374 -1843 91391 -1824
rect 88278 -3169 88302 -3142
rect 88283 -3403 88306 -3377
rect 93993 -1825 94015 -1800
rect 89707 -4826 89728 -4803
rect 89708 -4942 89729 -4919
rect 91381 -7426 91398 -7409
rect 91376 -7548 91393 -7531
<< metal1 >>
rect 97829 14454 97871 14461
rect 97829 14431 97841 14454
rect 97861 14431 97871 14454
rect 97829 14307 97871 14431
rect 97829 14284 97840 14307
rect 97860 14284 97871 14307
rect 97829 14274 97871 14284
rect 83075 2401 83119 2405
rect 83075 2384 83089 2401
rect 83108 2384 83119 2401
rect 83075 975 83119 2384
rect 83075 958 83087 975
rect 83106 958 83119 975
rect 83075 948 83119 958
rect 83399 977 83419 1557
rect 83399 922 83422 977
rect 83069 604 83103 606
rect 83069 600 83104 604
rect 83069 582 83075 600
rect 83092 582 83104 600
rect 83069 581 83104 582
rect 83070 579 83104 581
rect 83070 489 83093 579
rect 83401 511 83422 922
rect 86566 639 86611 667
rect 86566 612 86577 639
rect 86600 612 86611 639
rect 84887 597 84916 603
rect 84887 580 84893 597
rect 84910 580 84916 597
rect 84887 575 84916 580
rect 84889 516 84907 575
rect 83070 488 83073 489
rect 83069 470 83073 488
rect 83090 470 83093 489
rect 83394 501 83430 511
rect 83394 478 83402 501
rect 83424 478 83430 501
rect 84885 509 84914 516
rect 84885 492 84890 509
rect 84908 492 84914 509
rect 84885 486 84914 492
rect 83394 470 83430 478
rect 83069 462 83093 470
rect 86566 444 86611 612
rect 86566 417 86575 444
rect 86598 417 86611 444
rect 88274 623 88310 646
rect 88274 601 88284 623
rect 88302 601 88310 623
rect 88274 473 88310 601
rect 89701 615 89735 622
rect 89701 592 89707 615
rect 89728 592 89735 615
rect 89701 507 89735 592
rect 89701 484 89709 507
rect 89730 484 89735 507
rect 89701 474 89735 484
rect 91369 617 91394 628
rect 91369 598 91374 617
rect 91391 598 91394 617
rect 91369 475 91394 598
rect 88274 451 88284 473
rect 88302 451 88310 473
rect 88274 442 88310 451
rect 91369 456 91374 475
rect 91391 456 91394 475
rect 93988 623 94023 633
rect 93988 598 93996 623
rect 94018 598 94023 623
rect 93988 500 94023 598
rect 93988 475 93994 500
rect 94016 475 94023 500
rect 93988 467 94023 475
rect 91369 449 91394 456
rect 86566 403 86611 417
rect 101663 116 101710 119
rect 101663 88 101680 116
rect 101707 88 101710 116
rect 101663 82 101710 88
rect 102432 -47 102461 -37
rect 102432 -66 102435 -47
rect 102454 -66 102461 -47
rect 102432 -73 102461 -66
rect 101308 -270 101347 -249
rect 101308 -297 101314 -270
rect 101308 -298 101315 -297
rect 101341 -298 101347 -270
rect 101308 -315 101347 -298
rect 86565 -1384 86604 -1366
rect 89697 -1372 89729 -1344
rect 83279 -1420 83315 -1409
rect 83279 -1445 83284 -1420
rect 83306 -1445 83315 -1420
rect 86565 -1411 86575 -1384
rect 86598 -1411 86604 -1384
rect 83279 -1450 83315 -1445
rect 84811 -1433 84841 -1427
rect 83283 -2164 83297 -1450
rect 84811 -1454 84816 -1433
rect 84838 -1454 84841 -1433
rect 84811 -1459 84841 -1454
rect 84812 -1816 84839 -1459
rect 84808 -1824 84846 -1816
rect 84808 -1845 84814 -1824
rect 84836 -1845 84846 -1824
rect 84808 -1851 84846 -1845
rect 86565 -1840 86604 -1411
rect 86565 -1867 86576 -1840
rect 86599 -1867 86604 -1840
rect 86565 -1899 86604 -1867
rect 88274 -1385 88312 -1377
rect 88274 -1412 88281 -1385
rect 88305 -1412 88312 -1385
rect 88274 -1840 88312 -1412
rect 88274 -1867 88280 -1840
rect 88304 -1867 88312 -1840
rect 88274 -1875 88312 -1867
rect 89697 -1395 89704 -1372
rect 89725 -1395 89729 -1372
rect 89697 -1853 89729 -1395
rect 91371 -1402 91392 -1398
rect 91370 -1406 91394 -1402
rect 91369 -1407 91394 -1406
rect 91369 -1426 91373 -1407
rect 91390 -1426 91394 -1407
rect 95726 -1403 95766 -1385
rect 91369 -1428 91394 -1426
rect 93985 -1421 94024 -1413
rect 91369 -1432 91393 -1428
rect 91371 -1821 91392 -1432
rect 93985 -1446 93993 -1421
rect 94015 -1446 94024 -1421
rect 93985 -1800 94024 -1446
rect 95726 -1429 95736 -1403
rect 95760 -1429 95766 -1403
rect 95726 -1607 95766 -1429
rect 97830 -1428 97872 -1408
rect 97830 -1451 97843 -1428
rect 97864 -1451 97872 -1428
rect 97830 -1549 97872 -1451
rect 97830 -1572 97841 -1549
rect 97862 -1572 97872 -1549
rect 97830 -1580 97872 -1572
rect 95726 -1633 95730 -1607
rect 95754 -1633 95766 -1607
rect 95726 -1642 95766 -1633
rect 91371 -1824 91396 -1821
rect 91371 -1843 91374 -1824
rect 91391 -1843 91396 -1824
rect 93985 -1825 93993 -1800
rect 94015 -1825 94024 -1800
rect 93985 -1833 94024 -1825
rect 91371 -1847 91396 -1843
rect 91371 -1852 91392 -1847
rect 89697 -1876 89704 -1853
rect 89725 -1876 89729 -1853
rect 89697 -1891 89729 -1876
rect 83283 -2226 83301 -2164
rect 83280 -2227 83303 -2226
rect 83275 -2230 83309 -2227
rect 83275 -2245 83283 -2230
rect 83276 -2247 83283 -2245
rect 83301 -2247 83309 -2230
rect 83276 -2253 83309 -2247
rect 84809 -2375 84839 -2368
rect 84809 -2394 84817 -2375
rect 84835 -2394 84839 -2375
rect 84809 -2397 84839 -2394
rect 84812 -2471 84838 -2397
rect 84812 -2472 84842 -2471
rect 84811 -2476 84842 -2472
rect 84811 -2496 84816 -2476
rect 84837 -2496 84842 -2476
rect 84811 -2503 84842 -2496
rect 86564 -2802 86602 -2595
rect 88273 -3142 88311 -3123
rect 88273 -3169 88278 -3142
rect 88302 -3169 88311 -3142
rect 88273 -3365 88311 -3169
rect 88273 -3377 88313 -3365
rect 88273 -3403 88283 -3377
rect 88306 -3403 88313 -3377
rect 88273 -3408 88313 -3403
rect 88274 -3410 88313 -3408
rect 89700 -4803 89734 -4795
rect 89700 -4826 89707 -4803
rect 89728 -4826 89734 -4803
rect 89700 -4915 89734 -4826
rect 89700 -4919 89735 -4915
rect 89700 -4942 89708 -4919
rect 89729 -4942 89735 -4919
rect 89700 -4948 89735 -4942
rect 91375 -7409 91405 -7402
rect 91374 -7426 91381 -7409
rect 91398 -7426 91405 -7409
rect 91374 -7431 91405 -7426
rect 91374 -7525 91400 -7431
rect 91371 -7531 91401 -7525
rect 91371 -7548 91376 -7531
rect 91393 -7548 91401 -7531
rect 91371 -7554 91401 -7548
<< via1 >>
rect 101680 88 101707 116
rect 101314 -297 101341 -270
rect 101315 -298 101341 -297
<< metal2 >>
rect 98054 14085 98097 14469
rect 98054 13822 98099 14085
rect 83944 -1059 84003 -1054
rect 98060 -1059 98099 13822
rect 101675 161 101716 166
rect 101674 159 101716 161
rect 101674 128 101680 159
rect 101711 128 101716 159
rect 101674 121 101716 128
rect 101674 116 101710 121
rect 101674 88 101680 116
rect 101707 88 101710 116
rect 101674 82 101710 88
rect 101248 -265 101278 -261
rect 101248 -270 101344 -265
rect 101248 -297 101314 -270
rect 101248 -298 101315 -297
rect 101341 -298 101344 -270
rect 101248 -300 101344 -298
rect 101248 -1059 101278 -300
rect 83944 -1099 101278 -1059
rect 83944 -1907 84003 -1099
rect 98060 -1110 98099 -1099
<< via2 >>
rect 101680 128 101711 159
<< metal3 >>
rect 101673 218 101711 234
rect 101673 189 101677 218
rect 101674 185 101677 189
rect 101709 212 101711 218
rect 101709 185 101715 212
rect 101674 168 101715 185
rect 101675 159 101715 168
rect 101675 128 101680 159
rect 101711 128 101715 159
rect 101675 121 101715 128
<< via3 >>
rect 101677 185 101709 218
<< metal4 >>
rect 100581 15522 100759 15525
rect 98527 15489 100820 15522
rect 100581 15484 100820 15489
rect 100770 12714 100820 15484
rect 100770 12610 100867 12714
rect 100771 324 100867 12610
rect 100771 288 101710 324
rect 100777 207 100860 288
rect 101674 258 101710 288
rect 101673 248 101710 258
rect 101673 218 101711 248
rect 100777 157 100862 207
rect 101673 185 101677 218
rect 101709 212 101711 218
rect 101709 185 101717 212
rect 101673 176 101717 185
rect 83467 -814 83701 -812
rect 100779 -814 100862 157
rect 83467 -914 100862 -814
rect 83473 -1421 83532 -914
rect 83468 -1456 83532 -1421
rect 83468 -2006 83527 -1456
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 82880 0 1 2634
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 101227 0 1 -409
box 20 86 1230 590
use 9bitdac_layout  9bitdac_layout_1
timestamp 1616555653
transform 1 0 -214 0 1 -27858
box 0 -988 99386 26397
use 9bitdac_layout  9bitdac_layout_0
timestamp 1616555653
transform 1 0 0 0 1 988
box 0 -988 99386 26397
<< labels >>
rlabel locali 83001 2598 83001 2598 1 x1_vref5
rlabel locali 83089 2429 83089 2429 1 x2_vref1
rlabel locali 82797 -26253 82797 -26253 1 inp2
rlabel locali 415 26984 415 26984 1 inp1
rlabel locali 101212 -140 101212 -140 1 d9
rlabel locali 102481 -59 102481 -59 1 out_v
rlabel metal2 101269 -283 101269 -283 1 gnd!
rlabel metal4 101688 244 101688 244 1 vdd!
rlabel locali 102354 216 102354 216 1 x1_out_v
rlabel locali 102365 -356 102365 -356 1 x2_out_v
rlabel locali 83290 207 83290 207 1 d0
rlabel locali 84821 72 84821 72 1 d1
rlabel locali 86585 -283 86585 -283 1 d2
rlabel locali 88291 -430 88291 -430 1 d3
rlabel locali 89716 -172 89716 -172 1 d4
rlabel locali 91382 -85 91382 -85 1 d5
rlabel locali 94000 -69 94000 -69 1 d6
rlabel locali 95750 -475 95750 -475 1 d7
rlabel locali 97853 -610 97853 -610 1 d8
<< end >>
