* SPICE3 file created from 10bitdac_layout.ext - technology: sky130A

*Model Description
.para temp =27 

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 switch_layout_0/dd switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1 switch_layout_0/dd switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2 switch_layout_0/dinb d9 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3 switch_layout_0/dinb d9 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4 x1_out_v switch_layout_0/dd out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5 out_v switch_layout_0/dinb x1_out_v switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6 x2_out_v switch_layout_0/dd out_v switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7 out_v switch_layout_0/dinb x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8 x1_vref5 x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9 9bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X10 9bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X11 9bitdac_layout_0/switch_layout_0/dinb d8 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X12 9bitdac_layout_0/switch_layout_0/dinb d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X13 9bitdac_layout_0/x1_out_v 9bitdac_layout_0/switch_layout_0/dd x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X14 x1_out_v 9bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/x1_out_v 9bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X15 9bitdac_layout_0/x2_out_v 9bitdac_layout_0/switch_layout_0/dd x1_out_v 9bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X16 x1_out_v 9bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X17 9bitdac_layout_0/x1_vref5 9bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X18 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X19 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X20 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb d7 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X21 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X22 9bitdac_layout_0/8bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X23 9bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X24 9bitdac_layout_0/8bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X25 9bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X26 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X27 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X28 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X29 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X30 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X31 9bitdac_layout_0/8bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X32 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X33 9bitdac_layout_0/8bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X34 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X35 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X36 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X37 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X38 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X39 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X40 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X41 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X42 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X43 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X44 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X45 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X46 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X47 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X48 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X49 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X50 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X51 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X52 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X53 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X54 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X55 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X56 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X57 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X58 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X59 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X60 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X61 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X62 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X63 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X64 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X65 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X66 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X67 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X68 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X69 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X70 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X71 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X72 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X73 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X74 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X75 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X76 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X77 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X78 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X79 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X80 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X81 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X82 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X83 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X84 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X85 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X86 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X87 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X88 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X89 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X90 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X91 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X92 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X93 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X94 inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X95 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X96 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X97 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X98 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X99 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X100 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X101 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X102 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X103 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X104 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X105 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X106 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X107 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X108 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X109 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X110 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X111 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X112 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X113 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X114 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X115 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X116 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X117 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X118 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X119 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X120 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X121 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X122 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X123 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X124 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X125 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X126 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X127 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X128 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X129 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X130 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X131 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X132 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X133 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X134 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X135 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X136 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X137 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X138 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X139 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X140 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X141 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X142 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X143 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X144 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X145 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X146 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X147 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X148 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X149 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X150 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X151 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X152 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X153 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X154 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X155 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X156 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X157 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X158 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X159 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X160 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X161 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X162 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X163 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X164 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X165 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X166 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X167 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X168 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X169 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X170 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X171 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X172 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X173 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X174 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X175 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X176 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X177 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X178 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X179 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X180 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X181 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X182 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X183 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X184 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X185 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X186 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X187 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X188 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X189 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X190 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X191 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X192 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X193 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X194 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X195 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X196 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X197 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X198 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X199 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X200 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X201 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X202 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X203 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X204 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X205 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X206 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X207 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X208 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X209 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X210 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X211 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X212 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X213 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X214 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X215 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X216 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X217 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X218 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X219 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X220 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X221 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X222 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X223 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X224 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X225 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X226 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X227 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X228 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X229 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X230 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X231 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X232 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X233 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X234 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X235 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X236 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X237 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X238 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X239 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X240 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X241 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X242 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X243 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X244 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X245 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X246 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X247 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X248 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X249 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X250 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X251 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X252 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X253 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X254 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X255 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X256 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X257 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X258 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X259 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X260 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X261 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X262 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X263 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X264 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X265 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X266 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X267 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X268 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X269 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X270 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X271 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X272 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X273 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X274 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X275 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X276 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X277 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X278 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X279 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X280 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X281 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X282 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X283 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X284 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X285 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X286 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X287 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X288 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X289 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X290 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X291 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X292 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X293 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X294 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X295 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X296 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X297 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X298 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X299 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X300 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X301 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X302 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X303 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X304 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X305 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X306 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X307 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X308 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X309 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X310 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X311 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X312 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X313 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X314 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X315 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X316 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X317 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X318 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X319 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X320 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X321 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X322 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X323 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X324 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X325 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X326 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X327 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X328 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X329 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X330 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X331 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X332 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X333 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X334 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X335 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X336 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X337 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X338 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X339 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X340 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X341 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X342 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X343 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X344 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X345 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X346 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X347 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X348 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X349 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X350 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X351 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X352 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X353 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X354 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X355 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X356 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X357 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X358 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X359 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X360 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X361 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X362 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X363 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X364 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X365 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X366 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X367 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X368 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X369 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X370 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X371 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X372 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X373 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X374 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X375 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X376 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X377 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X378 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X379 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X380 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X381 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X382 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X383 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X384 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X385 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X386 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X387 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X388 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X389 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X390 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X391 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X392 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X393 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X394 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X395 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X396 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X397 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X398 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X399 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X400 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X401 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X402 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X403 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X404 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X405 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X406 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X407 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X408 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X409 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X410 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X411 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X412 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X413 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X414 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X415 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X416 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X417 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X418 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X419 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X420 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X421 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X422 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X423 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X424 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X425 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X426 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X427 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X428 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X429 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X430 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X431 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X432 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X433 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X434 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X435 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X436 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X437 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X438 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X439 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X440 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X441 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X442 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X443 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X444 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X445 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X446 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X447 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X448 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X449 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X450 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X451 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X452 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X453 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X454 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X455 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X456 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X457 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X458 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X459 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X460 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X461 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X462 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X463 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X464 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X465 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X466 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X467 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X468 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X469 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X470 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X471 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X472 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X473 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X474 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X475 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X476 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X477 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X478 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X479 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X480 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X481 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X482 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X483 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X484 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X485 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X486 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X487 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X488 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X489 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X490 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X491 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X492 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X493 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X494 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X495 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X496 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X497 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X498 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X499 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X500 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X501 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X502 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X503 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X504 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X505 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X506 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X507 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X508 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X509 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X510 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X511 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X512 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X513 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X514 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X515 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X516 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X517 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X518 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X519 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X520 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X521 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X522 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X523 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X524 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X525 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X526 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X527 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X528 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X529 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X530 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X531 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X532 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X533 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X534 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X535 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X536 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X537 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X538 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X539 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X540 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X541 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X542 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X543 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X544 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X545 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X546 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X547 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X548 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X549 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X550 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X551 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X552 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X553 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X554 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X555 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X556 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X557 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X558 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X559 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X560 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X561 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X562 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X563 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X564 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X565 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X566 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X567 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X568 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X569 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X570 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X571 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X572 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X573 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X574 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X575 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X576 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X577 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X578 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X579 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X580 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X581 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X582 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X583 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X584 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X585 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X586 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X587 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X588 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X589 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X590 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X591 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X592 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X593 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X594 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X595 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X596 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X597 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X598 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X599 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X600 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X601 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X602 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X603 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X604 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X605 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X606 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X607 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X608 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X609 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X610 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X611 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X612 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X613 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X614 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X615 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X616 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X617 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X618 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X619 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X620 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X621 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X622 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X623 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X624 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X625 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X626 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X627 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X628 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X629 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X630 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X631 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X632 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X633 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X634 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X635 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X636 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X637 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X638 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X639 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X640 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X641 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X642 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X643 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X644 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X645 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X646 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X647 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X648 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X649 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X650 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X651 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X652 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X653 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X654 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X655 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X656 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X657 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X658 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X659 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X660 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X661 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X662 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X663 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X664 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X665 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X666 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X667 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X668 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X669 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X670 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X671 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X672 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X673 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X674 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X675 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X676 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X677 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X678 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X679 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X680 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X681 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X682 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X683 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X684 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X685 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X686 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X687 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X688 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X689 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X690 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X691 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X692 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X693 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X694 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X695 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X696 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X697 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X698 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X699 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X700 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X701 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X702 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X703 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X704 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X705 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X706 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X707 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X708 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X709 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X710 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X711 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X712 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X713 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X714 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X715 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X716 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X717 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X718 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X719 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X720 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X721 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X722 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X723 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X724 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X725 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X726 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X727 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X728 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X729 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X730 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X731 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X732 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X733 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X734 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X735 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X736 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X737 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X738 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X739 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X740 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X741 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X742 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X743 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X744 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X745 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X746 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X747 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X748 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X749 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X750 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X751 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X752 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X753 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X754 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X755 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X756 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X757 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X758 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X759 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X760 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X761 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X762 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X763 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X764 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X765 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X766 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X767 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X768 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X769 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X770 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X771 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X772 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X773 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X774 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X775 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X776 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X777 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X778 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X779 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X780 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X781 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X782 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X783 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X784 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X785 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X786 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X787 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X788 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X789 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X790 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X791 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X792 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X793 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X794 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X795 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X796 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X797 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X798 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X799 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X800 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X801 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X802 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X803 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X804 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X805 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X806 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X807 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X808 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X809 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X810 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X811 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X812 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X813 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X814 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X815 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X816 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X817 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X818 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X819 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X820 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X821 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X822 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X823 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X824 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X825 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X826 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X827 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X828 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X829 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X830 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X831 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X832 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X833 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X834 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X835 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X836 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X837 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X838 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X839 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X840 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X841 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X842 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X843 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X844 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X845 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X846 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X847 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X848 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X849 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X850 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X851 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X852 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X853 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X854 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X855 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X856 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X857 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X858 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X859 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X860 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X861 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X862 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X863 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X864 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X865 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X866 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X867 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X868 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X869 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X870 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X871 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X872 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X873 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X874 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X875 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X876 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X877 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X878 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X879 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X880 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X881 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X882 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X883 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X884 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X885 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X886 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X887 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X888 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X889 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X890 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X891 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X892 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X893 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X894 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X895 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X896 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X897 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X898 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X899 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X900 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X901 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X902 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X903 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X904 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X905 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X906 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X907 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X908 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X909 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X910 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X911 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X912 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X913 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X914 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X915 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X916 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X917 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X918 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X919 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X920 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X921 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X922 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X923 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X924 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X925 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X926 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X927 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X928 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X929 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X930 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X931 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X932 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X933 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X934 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X935 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X936 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X937 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X938 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X939 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X940 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X941 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X942 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X943 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X944 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X945 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X946 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X947 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X948 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X949 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X950 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X951 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X952 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X953 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X954 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X955 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X956 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X957 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X958 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X959 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X960 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X961 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X962 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X963 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X964 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X965 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X966 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X967 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X968 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X969 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X970 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X971 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X972 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X973 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X974 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X975 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X976 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X977 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X978 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X979 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X980 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X981 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X982 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X983 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X984 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X985 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X986 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X987 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X988 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X989 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X990 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X991 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X992 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X993 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X994 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X995 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X996 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X997 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X998 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X999 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1000 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1001 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1002 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1003 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1004 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1005 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1006 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1007 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1008 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1009 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1010 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1011 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1012 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1013 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1014 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1015 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1016 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1017 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1018 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1019 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1020 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1021 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1022 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1023 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1024 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1025 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1026 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1027 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1028 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1029 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1030 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1031 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1032 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1033 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1034 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1035 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1036 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1037 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1038 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1039 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1040 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1041 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1042 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1043 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1044 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1045 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1046 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1047 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1048 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1049 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1050 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1051 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1052 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1053 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1054 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1055 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1056 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1057 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1058 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1059 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1060 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1061 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1062 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1063 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1064 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1065 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1066 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1067 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1068 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1069 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1070 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1071 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1072 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1073 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1074 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1075 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1076 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1077 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1078 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1079 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1080 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1081 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1082 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1083 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1084 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1085 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1086 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1087 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1088 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1089 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1090 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1091 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1092 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1093 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1094 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1095 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1096 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1097 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1098 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1099 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1100 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1101 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1102 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1103 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1104 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1105 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1106 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1107 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1108 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1109 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1110 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1111 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1112 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1113 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1114 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1115 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1116 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1117 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1118 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1119 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1120 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1121 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1122 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1123 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1124 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1125 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1126 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1127 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1128 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1129 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1130 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1131 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1132 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1133 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1134 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1135 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1136 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1137 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1138 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1139 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1140 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1141 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1142 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1143 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1144 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1145 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1146 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1147 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1148 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1149 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1150 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1151 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1152 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1153 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1154 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1155 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1156 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1157 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1158 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1159 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1160 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1161 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1162 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1163 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1164 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1165 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1166 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1167 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1168 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1169 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1170 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1171 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1172 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1173 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1174 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1175 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1176 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1177 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1178 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1179 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1180 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1181 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1182 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1183 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1184 9bitdac_layout_0/8bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1185 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1186 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1187 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1188 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1189 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1190 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1191 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1192 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1193 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1194 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1195 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1196 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1197 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1198 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1199 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1200 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1201 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1202 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1203 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1204 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1205 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1206 9bitdac_layout_0/8bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1207 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1208 9bitdac_layout_0/8bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1209 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1210 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1211 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1212 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1213 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1214 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1215 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1216 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1217 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1218 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1219 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1220 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1221 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1222 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1223 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1224 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1225 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1226 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1227 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1228 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1229 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1230 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1231 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1232 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1233 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1234 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1235 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1236 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1237 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1238 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1239 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1240 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1241 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1242 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1243 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1244 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1245 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1246 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1247 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1248 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1249 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1250 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1251 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1252 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1253 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1254 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1255 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1256 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1257 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1258 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1259 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1260 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1261 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1262 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1263 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1264 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1265 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1266 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1267 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1268 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1269 9bitdac_layout_0/8bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1270 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1271 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1272 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1273 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1274 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1275 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1276 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1277 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1278 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1279 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1280 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1281 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1282 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1283 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1284 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1285 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1286 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1287 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1288 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1289 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1290 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1291 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1292 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1293 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1294 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1295 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1296 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1297 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1298 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1299 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1300 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1301 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1302 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1303 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1304 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1305 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1306 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1307 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1308 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1309 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1310 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1311 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1312 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1313 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1314 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1315 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1316 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1317 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1318 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1319 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1320 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1321 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1322 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1323 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1324 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1325 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1326 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1327 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1328 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1329 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1330 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1331 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1332 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1333 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1334 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1335 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1336 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1337 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1338 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1339 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1340 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1341 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1342 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1343 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1344 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1345 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1346 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1347 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1348 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1349 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1350 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1351 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1352 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1353 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1354 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1355 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1356 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1357 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1358 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1359 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1360 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1361 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1362 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1363 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1364 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1365 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1366 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1367 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1368 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1369 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1370 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1371 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1372 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1373 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1374 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1375 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1376 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1377 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1378 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1379 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1380 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1381 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1382 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1383 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1384 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1385 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1386 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1387 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1388 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1389 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1390 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1391 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1392 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1393 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1394 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1395 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1396 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1397 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1398 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1399 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1400 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1401 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1402 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1403 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1404 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1405 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1406 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1407 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1408 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1409 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1410 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1411 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1412 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1413 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1414 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1415 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1416 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1417 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1418 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1419 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1420 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1421 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1422 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1423 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1424 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1425 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1426 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1427 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1428 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1429 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1430 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1431 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1432 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1433 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1434 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1435 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1436 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1437 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1438 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1439 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1440 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1441 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1442 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1443 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1444 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1445 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1446 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1447 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1448 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1449 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1450 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1451 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1452 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1453 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1454 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1455 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1456 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1457 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1458 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1459 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1460 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1461 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1462 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1463 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1464 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1465 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1466 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1467 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1468 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1469 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1470 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1471 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1472 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1473 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1474 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1475 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1476 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1477 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1478 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1479 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1480 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1481 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1482 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1483 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1484 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1485 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1486 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1487 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1488 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1489 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1490 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1491 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1492 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1493 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1494 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1495 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1496 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1497 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1498 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1499 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1500 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1501 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1502 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1503 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1504 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1505 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1506 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1507 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1508 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1509 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1510 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1511 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1512 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1513 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1514 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1515 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1516 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1517 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1518 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1519 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1520 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1521 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1522 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1523 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1524 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1525 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1526 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1527 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1528 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1529 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1530 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1531 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1532 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1533 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1534 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1535 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1536 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1537 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1538 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1539 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1540 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1541 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1542 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1543 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1544 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1545 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1546 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1547 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1548 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1549 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1550 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1551 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1552 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1553 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1554 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1555 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1556 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1557 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1558 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1559 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1560 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1561 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1562 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1563 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1564 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1565 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1566 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1567 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1568 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1569 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1570 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1571 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1572 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1573 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1574 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1575 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1576 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1577 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1578 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1579 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1580 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1581 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1582 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1583 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1584 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1585 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1586 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1587 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1588 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1589 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1590 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1591 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1592 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1593 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1594 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1595 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1596 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1597 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1598 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1599 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1600 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1601 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1602 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1603 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1604 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1605 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1606 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1607 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1608 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1609 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1610 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1611 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1612 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1613 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1614 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1615 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1616 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1617 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1618 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1619 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1620 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1621 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1622 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1623 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1624 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1625 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1626 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1627 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1628 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1629 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1630 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1631 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1632 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1633 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1634 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1635 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1636 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1637 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1638 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1639 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1640 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1641 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1642 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1643 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1644 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1645 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1646 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1647 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1648 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1649 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1650 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1651 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1652 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1653 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1654 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1655 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1656 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1657 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1658 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1659 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1660 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1661 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1662 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1663 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1664 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1665 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1666 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1667 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1668 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1669 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1670 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1671 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1672 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1673 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1674 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1675 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1676 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1677 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1678 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1679 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1680 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1681 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1682 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1683 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1684 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1685 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1686 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1687 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1688 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1689 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1690 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1691 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1692 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1693 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1694 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1695 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1696 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1697 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1698 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1699 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1700 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1701 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1702 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1703 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1704 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1705 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1706 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1707 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1708 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1709 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1710 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1711 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1712 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1713 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1714 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1715 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1716 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1717 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1718 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1719 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1720 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1721 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1722 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1723 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1724 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1725 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1726 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1727 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1728 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1729 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1730 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1731 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1732 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1733 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1734 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1735 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1736 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1737 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1738 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1739 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1740 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1741 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1742 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1743 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1744 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1745 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1746 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1747 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1748 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1749 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1750 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1751 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1752 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1753 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1754 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1755 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1756 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1757 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1758 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1759 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1760 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1761 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1762 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1763 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1764 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1765 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1766 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1767 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1768 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1769 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1770 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1771 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1772 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1773 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1774 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1775 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1776 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1777 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1778 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1779 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1780 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1781 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1782 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1783 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1784 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1785 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1786 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1787 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1788 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1789 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1790 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1791 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1792 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1793 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1794 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1795 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1796 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1797 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1798 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1799 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1800 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1801 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1802 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1803 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1804 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1805 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1806 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1807 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1808 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1809 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1810 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1811 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1812 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1813 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1814 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1815 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1816 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1817 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1818 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1819 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1820 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1821 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1822 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1823 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1824 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1825 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1826 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1827 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1828 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1829 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1830 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1831 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1832 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1833 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1834 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1835 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1836 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1837 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1838 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1839 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1840 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1841 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1842 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1843 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1844 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1845 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1846 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1847 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1848 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1849 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1850 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1851 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1852 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1853 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1854 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1855 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1856 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1857 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1858 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1859 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1860 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1861 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1862 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1863 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1864 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1865 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1866 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1867 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1868 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1869 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1870 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1871 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1872 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1873 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1874 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1875 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1876 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1877 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1878 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1879 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1880 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1881 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1882 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1883 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1884 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1885 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1886 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1887 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1888 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1889 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1890 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1891 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1892 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1893 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1894 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1895 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1896 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1897 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1898 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1899 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1900 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1901 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1902 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1903 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1904 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1905 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1906 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1907 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1908 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1909 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1910 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1911 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1912 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1913 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1914 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1915 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1916 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1917 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1918 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1919 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1920 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1921 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1922 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1923 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1924 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1925 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1926 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1927 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1928 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1929 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1930 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1931 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1932 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1933 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1934 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1935 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1936 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1937 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1938 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1939 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1940 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1941 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1942 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1943 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1944 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1945 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1946 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1947 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1948 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1949 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1950 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1951 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1952 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1953 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1954 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1955 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1956 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1957 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1958 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1959 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1960 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1961 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1962 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1963 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1964 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1965 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1966 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1967 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1968 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1969 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1970 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1971 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1972 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1973 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1974 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1975 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1976 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1977 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1978 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1979 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1980 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1981 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1982 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1983 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1984 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1985 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1986 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1987 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1988 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1989 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1990 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1991 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X1992 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X1993 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1994 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1995 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X1996 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X1997 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X1998 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X1999 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2000 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2001 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2002 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2003 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2004 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2005 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2006 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2007 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2008 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2009 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2010 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2011 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2012 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2013 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2014 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2015 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2016 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2017 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2018 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2019 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2020 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2021 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2022 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2023 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2024 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2025 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2026 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2027 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2028 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2029 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2030 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2031 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2032 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2033 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2034 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2035 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2036 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2037 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2038 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2039 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2040 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2041 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2042 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2043 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2044 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2045 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2046 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2047 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2048 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2049 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2050 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2051 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2052 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2053 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2054 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2055 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2056 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2057 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2058 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2059 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2060 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2061 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2062 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2063 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2064 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2065 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2066 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2067 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2068 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2069 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2070 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2071 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2072 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2073 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2074 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2075 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2076 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2077 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2078 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2079 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2080 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2081 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2082 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2083 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2084 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2085 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2086 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2087 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2088 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2089 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2090 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2091 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2092 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2093 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2094 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2095 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2096 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2097 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2098 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2099 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2100 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2101 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2102 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2103 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2104 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2105 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2106 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2107 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2108 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2109 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2110 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2111 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2112 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2113 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2114 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2115 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2116 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2117 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2118 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2119 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2120 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2121 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2122 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2123 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2124 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2125 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2126 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2127 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2128 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2129 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2130 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2131 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2132 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2133 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2134 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2135 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2136 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2137 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2138 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2139 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2140 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2141 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2142 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2143 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2144 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2145 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2146 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2147 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2148 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2149 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2150 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2151 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2152 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2153 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2154 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2155 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2156 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2157 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2158 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2159 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2160 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2161 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2162 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2163 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2164 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2165 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2166 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2167 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2168 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2169 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2170 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2171 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2172 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2173 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2174 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2175 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2176 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2177 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2178 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2179 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2180 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2181 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2182 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2183 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2184 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2185 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2186 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2187 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2188 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2189 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2190 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2191 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2192 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2193 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2194 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2195 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2196 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2197 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2198 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2199 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2200 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2201 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2202 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2203 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2204 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2205 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2206 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2207 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2208 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2209 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2210 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2211 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2212 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2213 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2214 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2215 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2216 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2217 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2218 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2219 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2220 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2221 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2222 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2223 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2224 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2225 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2226 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2227 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2228 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2229 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2230 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2231 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2232 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2233 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2234 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2235 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2236 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2237 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2238 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2239 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2240 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2241 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2242 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2243 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2244 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2245 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2246 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2247 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2248 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2249 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2250 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2251 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2252 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2253 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2254 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2255 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2256 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2257 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2258 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2259 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2260 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2261 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2262 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2263 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2264 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2265 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2266 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2267 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2268 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2269 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2270 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2271 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2272 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2273 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2274 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2275 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2276 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2277 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2278 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2279 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2280 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2281 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2282 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2283 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2284 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2285 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2286 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2287 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2288 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2289 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2290 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2291 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2292 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2293 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2294 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2295 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2296 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2297 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2298 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2299 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2300 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2301 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2302 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2303 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2304 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2305 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2306 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2307 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2308 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2309 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2310 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2311 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2312 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2313 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2314 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2315 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2316 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2317 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2318 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2319 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2320 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2321 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2322 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2323 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2324 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2325 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2326 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2327 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2328 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2329 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2330 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2331 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2332 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2333 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2334 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2335 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2336 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2337 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2338 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2339 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2340 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2341 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2342 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2343 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2344 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2345 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2346 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2347 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2348 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2349 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2350 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2351 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2352 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2353 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2354 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2355 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2356 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2357 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2358 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2359 9bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2360 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2361 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2362 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2363 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2364 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2365 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2366 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2367 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2368 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2369 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2370 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2371 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2372 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2373 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2374 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2375 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2376 9bitdac_layout_0/8bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2377 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2378 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2379 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb d7 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2380 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2381 9bitdac_layout_0/8bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2382 9bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2383 9bitdac_layout_0/8bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2384 9bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2385 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2386 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2387 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2388 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2389 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2390 9bitdac_layout_0/8bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2391 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2392 9bitdac_layout_0/8bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2393 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2394 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2395 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2396 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2397 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2398 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2399 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2400 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2401 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2402 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2403 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2404 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2405 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2406 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2407 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2408 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2409 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2410 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2411 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2412 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2413 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2414 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2415 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2416 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2417 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2418 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2419 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2420 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2421 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2422 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2423 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2424 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2425 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2426 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2427 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2428 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2429 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2430 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2431 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2432 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2433 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2434 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2435 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2436 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2437 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2438 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2439 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2440 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2441 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2442 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2443 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2444 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2445 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2446 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2447 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2448 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2449 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2450 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2451 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2452 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2453 9bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2454 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2455 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2456 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2457 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2458 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2459 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2460 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2461 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2462 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2463 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2464 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2465 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2466 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2467 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2468 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2469 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2470 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2471 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2472 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2473 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2474 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2475 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2476 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2477 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2478 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2479 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2480 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2481 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2482 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2483 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2484 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2485 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2486 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2487 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2488 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2489 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2490 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2491 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2492 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2493 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2494 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2495 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2496 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2497 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2498 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2499 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2500 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2501 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2502 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2503 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2504 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2505 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2506 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2507 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2508 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2509 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2510 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2511 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2512 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2513 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2514 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2515 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2516 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2517 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2518 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2519 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2520 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2521 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2522 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2523 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2524 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2525 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2526 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2527 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2528 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2529 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2530 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2531 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2532 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2533 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2534 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2535 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2536 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2537 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2538 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2539 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2540 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2541 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2542 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2543 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2544 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2545 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2546 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2547 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2548 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2549 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2550 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2551 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2552 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2553 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2554 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2555 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2556 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2557 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2558 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2559 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2560 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2561 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2562 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2563 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2564 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2565 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2566 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2567 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2568 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2569 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2570 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2571 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2572 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2573 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2574 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2575 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2576 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2577 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2578 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2579 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2580 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2581 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2582 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2583 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2584 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2585 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2586 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2587 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2588 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2589 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2590 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2591 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2592 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2593 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2594 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2595 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2596 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2597 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2598 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2599 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2600 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2601 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2602 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2603 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2604 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2605 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2606 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2607 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2608 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2609 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2610 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2611 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2612 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2613 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2614 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2615 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2616 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2617 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2618 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2619 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2620 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2621 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2622 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2623 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2624 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2625 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2626 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2627 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2628 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2629 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2630 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2631 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2632 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2633 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2634 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2635 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2636 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2637 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2638 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2639 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2640 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2641 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2642 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2643 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2644 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2645 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2646 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2647 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2648 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2649 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2650 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2651 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2652 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2653 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2654 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2655 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2656 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2657 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2658 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2659 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2660 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2661 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2662 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2663 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2664 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2665 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2666 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2667 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2668 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2669 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2670 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2671 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2672 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2673 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2674 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2675 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2676 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2677 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2678 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2679 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2680 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2681 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2682 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2683 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2684 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2685 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2686 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2687 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2688 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2689 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2690 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2691 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2692 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2693 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2694 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2695 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2696 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2697 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2698 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2699 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2700 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2701 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2702 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2703 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2704 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2705 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2706 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2707 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2708 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2709 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2710 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2711 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2712 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2713 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2714 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2715 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2716 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2717 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2718 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2719 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2720 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2721 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2722 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2723 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2724 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2725 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2726 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2727 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2728 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2729 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2730 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2731 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2732 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2733 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2734 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2735 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2736 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2737 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2738 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2739 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2740 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2741 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2742 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2743 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2744 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2745 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2746 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2747 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2748 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2749 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2750 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2751 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2752 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2753 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2754 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2755 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2756 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2757 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2758 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2759 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2760 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2761 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2762 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2763 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2764 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2765 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2766 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2767 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2768 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2769 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2770 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2771 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2772 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2773 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2774 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2775 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2776 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2777 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2778 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2779 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2780 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2781 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2782 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2783 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2784 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2785 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2786 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2787 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2788 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2789 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2790 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2791 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2792 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2793 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2794 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2795 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2796 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2797 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2798 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2799 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2800 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2801 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2802 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2803 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2804 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2805 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2806 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2807 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2808 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2809 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2810 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2811 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2812 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2813 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2814 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2815 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2816 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2817 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2818 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2819 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2820 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2821 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2822 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2823 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2824 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2825 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2826 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2827 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2828 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2829 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2830 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2831 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2832 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2833 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2834 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2835 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2836 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2837 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2838 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2839 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2840 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2841 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2842 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2843 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2844 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2845 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2846 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2847 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2848 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2849 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2850 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2851 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2852 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2853 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2854 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2855 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2856 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2857 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2858 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2859 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2860 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2861 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2862 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2863 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2864 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2865 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2866 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2867 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2868 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2869 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2870 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2871 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2872 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2873 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2874 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2875 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2876 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2877 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2878 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2879 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2880 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2881 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2882 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2883 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2884 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2885 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2886 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2887 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2888 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2889 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2890 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2891 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2892 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2893 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2894 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2895 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2896 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2897 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2898 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2899 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2900 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2901 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2902 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2903 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2904 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2905 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2906 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2907 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2908 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2909 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2910 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2911 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2912 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2913 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2914 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2915 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2916 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2917 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2918 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2919 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2920 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2921 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2922 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2923 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2924 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2925 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2926 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2927 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2928 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2929 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2930 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2931 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2932 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2933 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2934 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2935 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2936 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2937 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2938 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2939 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2940 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2941 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2942 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2943 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2944 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2945 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2946 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2947 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2948 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2949 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2950 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2951 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2952 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2953 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2954 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2955 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2956 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2957 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2958 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2959 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2960 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2961 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2962 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2963 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2964 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2965 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2966 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2967 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2968 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2969 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2970 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2971 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2972 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X2973 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2974 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2975 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2976 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2977 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2978 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2979 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2980 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2981 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2982 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2983 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2984 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2985 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2986 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2987 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2988 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2989 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2990 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X2991 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2992 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2993 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X2994 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2995 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2996 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X2997 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X2998 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X2999 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3000 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3001 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3002 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3003 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3004 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3005 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3006 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3007 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3008 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3009 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3010 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3011 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3012 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3013 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3014 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3015 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3016 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3017 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3018 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3019 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3020 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3021 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3022 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3023 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3024 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3025 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3026 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3027 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3028 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3029 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3030 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3031 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3032 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3033 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3034 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3035 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3036 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3037 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3038 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3039 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3040 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3041 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3042 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3043 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3044 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3045 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3046 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3047 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3048 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3049 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3050 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3051 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3052 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3053 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3054 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3055 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3056 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3057 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3058 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3059 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3060 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3061 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3062 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3063 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3064 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3065 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3066 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3067 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3068 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3069 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3070 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3071 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3072 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3073 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3074 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3075 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3076 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3077 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3078 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3079 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3080 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3081 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3082 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3083 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3084 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3085 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3086 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3087 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3088 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3089 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3090 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3091 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3092 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3093 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3094 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3095 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3096 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3097 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3098 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3099 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3100 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3101 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3102 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3103 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3104 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3105 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3106 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3107 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3108 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3109 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3110 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3111 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3112 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3113 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3114 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3115 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3116 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3117 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3118 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3119 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3120 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3121 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3122 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3123 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3124 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3125 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3126 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3127 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3128 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3129 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3130 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3131 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3132 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3133 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3134 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3135 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3136 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3137 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3138 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3139 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3140 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3141 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3142 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3143 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3144 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3145 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3146 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3147 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3148 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3149 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3150 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3151 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3152 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3153 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3154 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3155 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3156 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3157 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3158 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3159 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3160 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3161 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3162 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3163 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3164 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3165 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3166 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3167 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3168 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3169 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3170 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3171 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3172 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3173 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3174 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3175 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3176 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3177 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3178 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3179 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3180 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3181 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3182 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3183 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3184 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3185 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3186 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3187 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3188 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3189 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3190 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3191 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3192 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3193 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3194 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3195 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3196 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3197 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3198 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3199 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3200 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3201 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3202 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3203 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3204 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3205 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3206 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3207 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3208 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3209 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3210 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3211 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3212 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3213 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3214 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3215 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3216 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3217 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3218 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3219 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3220 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3221 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3222 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3223 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3224 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3225 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3226 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3227 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3228 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3229 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3230 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3231 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3232 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3233 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3234 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3235 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3236 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3237 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3238 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3239 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3240 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3241 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3242 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3243 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3244 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3245 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3246 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3247 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3248 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3249 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3250 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3251 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3252 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3253 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3254 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3255 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3256 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3257 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3258 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3259 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3260 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3261 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3262 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3263 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3264 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3265 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3266 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3267 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3268 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3269 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3270 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3271 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3272 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3273 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3274 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3275 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3276 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3277 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3278 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3279 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3280 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3281 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3282 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3283 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3284 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3285 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3286 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3287 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3288 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3289 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3290 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3291 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3292 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3293 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3294 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3295 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3296 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3297 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3298 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3299 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3300 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3301 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3302 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3303 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3304 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3305 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3306 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3307 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3308 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3309 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3310 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3311 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3312 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3313 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3314 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3315 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3316 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3317 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3318 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3319 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3320 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3321 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3322 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3323 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3324 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3325 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3326 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3327 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3328 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3329 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3330 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3331 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3332 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3333 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3334 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3335 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3336 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3337 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3338 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3339 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3340 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3341 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3342 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3343 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3344 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3345 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3346 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3347 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3348 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3349 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3350 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3351 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3352 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3353 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3354 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3355 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3356 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3357 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3358 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3359 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3360 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3361 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3362 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3363 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3364 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3365 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3366 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3367 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3368 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3369 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3370 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3371 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3372 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3373 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3374 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3375 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3376 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3377 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3378 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3379 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3380 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3381 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3382 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3383 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3384 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3385 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3386 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3387 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3388 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3389 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3390 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3391 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3392 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3393 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3394 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3395 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3396 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3397 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3398 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3399 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3400 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3401 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3402 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3403 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3404 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3405 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3406 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3407 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3408 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3409 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3410 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3411 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3412 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3413 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3414 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3415 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3416 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3417 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3418 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3419 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3420 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3421 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3422 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3423 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3424 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3425 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3426 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3427 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3428 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3429 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3430 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3431 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3432 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3433 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3434 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3435 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3436 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3437 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3438 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3439 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3440 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3441 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3442 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3443 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3444 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3445 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3446 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3447 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3448 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3449 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3450 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3451 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3452 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3453 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3454 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3455 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3456 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3457 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3458 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3459 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3460 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3461 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3462 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3463 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3464 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3465 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3466 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3467 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3468 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3469 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3470 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3471 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3472 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3473 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3474 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3475 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3476 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3477 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3478 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3479 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3480 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3481 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3482 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3483 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3484 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3485 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3486 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3487 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3488 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3489 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3490 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3491 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3492 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3493 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3494 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3495 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3496 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3497 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3498 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3499 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3500 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3501 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3502 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3503 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3504 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3505 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3506 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3507 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3508 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3509 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3510 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3511 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3512 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3513 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3514 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3515 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3516 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3517 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3518 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3519 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3520 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3521 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3522 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3523 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3524 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3525 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3526 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3527 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3528 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3529 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3530 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3531 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3532 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3533 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3534 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3535 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3536 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3537 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3538 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3539 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3540 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3541 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3542 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3543 9bitdac_layout_0/8bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3544 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3545 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3546 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3547 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3548 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3549 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3550 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3551 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3552 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3553 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3554 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3555 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3556 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3557 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3558 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3559 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3560 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3561 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3562 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3563 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3564 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3565 9bitdac_layout_0/8bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3566 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3567 9bitdac_layout_0/8bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3568 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3569 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3570 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3571 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3572 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3573 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3574 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3575 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3576 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3577 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3578 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3579 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3580 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3581 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3582 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3583 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3584 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3585 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3586 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3587 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3588 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3589 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3590 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3591 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3592 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3593 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3594 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3595 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3596 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3597 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3598 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3599 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3600 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3601 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3602 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3603 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3604 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3605 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3606 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3607 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3608 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3609 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3610 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3611 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3612 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3613 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3614 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3615 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3616 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3617 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3618 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3619 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3620 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3621 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3622 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3623 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3624 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3625 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3626 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3627 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3628 9bitdac_layout_0/8bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3629 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3630 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3631 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3632 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3633 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3634 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3635 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3636 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3637 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3638 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3639 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3640 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3641 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3642 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3643 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3644 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3645 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3646 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3647 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3648 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3649 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3650 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3651 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3652 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3653 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3654 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3655 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3656 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3657 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3658 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3659 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3660 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3661 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3662 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3663 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3664 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3665 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3666 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3667 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3668 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3669 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3670 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3671 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3672 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3673 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3674 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3675 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3676 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3677 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3678 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3679 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3680 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3681 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3682 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3683 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3684 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3685 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3686 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3687 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3688 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3689 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3690 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3691 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3692 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3693 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3694 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3695 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3696 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3697 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3698 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3699 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3700 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3701 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3702 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3703 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3704 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3705 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3706 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3707 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3708 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3709 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3710 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3711 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3712 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3713 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3714 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3715 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3716 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3717 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3718 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3719 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3720 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3721 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3722 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3723 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3724 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3725 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3726 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3727 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3728 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3729 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3730 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3731 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3732 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3733 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3734 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3735 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3736 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3737 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3738 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3739 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3740 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3741 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3742 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3743 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3744 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3745 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3746 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3747 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3748 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3749 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3750 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3751 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3752 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3753 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3754 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3755 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3756 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3757 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3758 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3759 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3760 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3761 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3762 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3763 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3764 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3765 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3766 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3767 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3768 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3769 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3770 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3771 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3772 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3773 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3774 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3775 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3776 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3777 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3778 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3779 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3780 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3781 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3782 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3783 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3784 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3785 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3786 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3787 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3788 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3789 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3790 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3791 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3792 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3793 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3794 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3795 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3796 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3797 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3798 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3799 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3800 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3801 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3802 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3803 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3804 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3805 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3806 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3807 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3808 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3809 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3810 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3811 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3812 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3813 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3814 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3815 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3816 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3817 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3818 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3819 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3820 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3821 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3822 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3823 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3824 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3825 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3826 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3827 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3828 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3829 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3830 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3831 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3832 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3833 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3834 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3835 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3836 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3837 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3838 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3839 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3840 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3841 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3842 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3843 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3844 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3845 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3846 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3847 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3848 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3849 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3850 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3851 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3852 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3853 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3854 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3855 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3856 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3857 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3858 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3859 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3860 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3861 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3862 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3863 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3864 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3865 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3866 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3867 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3868 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3869 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3870 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3871 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3872 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3873 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3874 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3875 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3876 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3877 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3878 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3879 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3880 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3881 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3882 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3883 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3884 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3885 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3886 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3887 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3888 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3889 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3890 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3891 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3892 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3893 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3894 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3895 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3896 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3897 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3898 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3899 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3900 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3901 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3902 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3903 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3904 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3905 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3906 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3907 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3908 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3909 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3910 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3911 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3912 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3913 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3914 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3915 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3916 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3917 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3918 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3919 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3920 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3921 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3922 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3923 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3924 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3925 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3926 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3927 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3928 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3929 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3930 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3931 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3932 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3933 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3934 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3935 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3936 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3937 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3938 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3939 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3940 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3941 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3942 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3943 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3944 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3945 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3946 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3947 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3948 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3949 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3950 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3951 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3952 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3953 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3954 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3955 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3956 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3957 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3958 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3959 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3960 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3961 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3962 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3963 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3964 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3965 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3966 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3967 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3968 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3969 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3970 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3971 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3972 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3973 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3974 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3975 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3976 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3977 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3978 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3979 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3980 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X3981 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X3982 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3983 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3984 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3985 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3986 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3987 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3988 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3989 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3990 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3991 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3992 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3993 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3994 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3995 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X3996 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X3997 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X3998 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X3999 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4000 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4001 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4002 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4003 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4004 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4005 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4006 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4007 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4008 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4009 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4010 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4011 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4012 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4013 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4014 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4015 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4016 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4017 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4018 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4019 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4020 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4021 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4022 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4023 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4024 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4025 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4026 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4027 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4028 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4029 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4030 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4031 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4032 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4033 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4034 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4035 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4036 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4037 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4038 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4039 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4040 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4041 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4042 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4043 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4044 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4045 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4046 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4047 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4048 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4049 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4050 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4051 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4052 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4053 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4054 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4055 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4056 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4057 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4058 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4059 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4060 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4061 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4062 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4063 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4064 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4065 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4066 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4067 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4068 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4069 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4070 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4071 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4072 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4073 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4074 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4075 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4076 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4077 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4078 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4079 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4080 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4081 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4082 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4083 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4084 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4085 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4086 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4087 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4088 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4089 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4090 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4091 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4092 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4093 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4094 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4095 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4096 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4097 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4098 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4099 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4100 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4101 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4102 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4103 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4104 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4105 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4106 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4107 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4108 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4109 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4110 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4111 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4112 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4113 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4114 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4115 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4116 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4117 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4118 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4119 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4120 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4121 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4122 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4123 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4124 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4125 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4126 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4127 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4128 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4129 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4130 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4131 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4132 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4133 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4134 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4135 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4136 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4137 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4138 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4139 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4140 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4141 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4142 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4143 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4144 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4145 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4146 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4147 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4148 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4149 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4150 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4151 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4152 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4153 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4154 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4155 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4156 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4157 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4158 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4159 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4160 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4161 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4162 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4163 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4164 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4165 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4166 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4167 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4168 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4169 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4170 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4171 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4172 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4173 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4174 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4175 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4176 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4177 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4178 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4179 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4180 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4181 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4182 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4183 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4184 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4185 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4186 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4187 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4188 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4189 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4190 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4191 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4192 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4193 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4194 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4195 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4196 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4197 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4198 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4199 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4200 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4201 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4202 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4203 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4204 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4205 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4206 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4207 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4208 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4209 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4210 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4211 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4212 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4213 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4214 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4215 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4216 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4217 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4218 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4219 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4220 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4221 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4222 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4223 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4224 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4225 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4226 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4227 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4228 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4229 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4230 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4231 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4232 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4233 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4234 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4235 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4236 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4237 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4238 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4239 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4240 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4241 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4242 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4243 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4244 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4245 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4246 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4247 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4248 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4249 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4250 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4251 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4252 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4253 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4254 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4255 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4256 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4257 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4258 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4259 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4260 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4261 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4262 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4263 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4264 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4265 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4266 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4267 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4268 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4269 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4270 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4271 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4272 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4273 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4274 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4275 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4276 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4277 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4278 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4279 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4280 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4281 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4282 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4283 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4284 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4285 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4286 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4287 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4288 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4289 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4290 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4291 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4292 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4293 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4294 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4295 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4296 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4297 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4298 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4299 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4300 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4301 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4302 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4303 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4304 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4305 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4306 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4307 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4308 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4309 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4310 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4311 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4312 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4313 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4314 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4315 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4316 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4317 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4318 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4319 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4320 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4321 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4322 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4323 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4324 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4325 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4326 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4327 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4328 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4329 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4330 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4331 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4332 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4333 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4334 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4335 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4336 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4337 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4338 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4339 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4340 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4341 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4342 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4343 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4344 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4345 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4346 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4347 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4348 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4349 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4350 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4351 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4352 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4353 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4354 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4355 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4356 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4357 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4358 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4359 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4360 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4361 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4362 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4363 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4364 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4365 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4366 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4367 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4368 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4369 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4370 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4371 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4372 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4373 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4374 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4375 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4376 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4377 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4378 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4379 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4380 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4381 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4382 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4383 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4384 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4385 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4386 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4387 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4388 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4389 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4390 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4391 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4392 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4393 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4394 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4395 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4396 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4397 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4398 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4399 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4400 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4401 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4402 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4403 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4404 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4405 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4406 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4407 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4408 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4409 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4410 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4411 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4412 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4413 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4414 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4415 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4416 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4417 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4418 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4419 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4420 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4421 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4422 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4423 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4424 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4425 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4426 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4427 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4428 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4429 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4430 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4431 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4432 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4433 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4434 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4435 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4436 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4437 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4438 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4439 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4440 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4441 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4442 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4443 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4444 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4445 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4446 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4447 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4448 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4449 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4450 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4451 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4452 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4453 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4454 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4455 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4456 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4457 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4458 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4459 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4460 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4461 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4462 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4463 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4464 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4465 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4466 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4467 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4468 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4469 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4470 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4471 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4472 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4473 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4474 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4475 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4476 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4477 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4478 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4479 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4480 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4481 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4482 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4483 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4484 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4485 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4486 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4487 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4488 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4489 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4490 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4491 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4492 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4493 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4494 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4495 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4496 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4497 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4498 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4499 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4500 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4501 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4502 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4503 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4504 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4505 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4506 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4507 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4508 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4509 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4510 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4511 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4512 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4513 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4514 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4515 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4516 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4517 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4518 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4519 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4520 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4521 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4522 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4523 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4524 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4525 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4526 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4527 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4528 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4529 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4530 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4531 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4532 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4533 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4534 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4535 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4536 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4537 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4538 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4539 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4540 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4541 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4542 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4543 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4544 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4545 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4546 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4547 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4548 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4549 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4550 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4551 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4552 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4553 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4554 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4555 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4556 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4557 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4558 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4559 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4560 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4561 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4562 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4563 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4564 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4565 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4566 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4567 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4568 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4569 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4570 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4571 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4572 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4573 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4574 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4575 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4576 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4577 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4578 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4579 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4580 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4581 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4582 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4583 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4584 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4585 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4586 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4587 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4588 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4589 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4590 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4591 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4592 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4593 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4594 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4595 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4596 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4597 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4598 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4599 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4600 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4601 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4602 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4603 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4604 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4605 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4606 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4607 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4608 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4609 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4610 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4611 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4612 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4613 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4614 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4615 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4616 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4617 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4618 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4619 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4620 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4621 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4622 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4623 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4624 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4625 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4626 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4627 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4628 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4629 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4630 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4631 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4632 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4633 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4634 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4635 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4636 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4637 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4638 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4639 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4640 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4641 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4642 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4643 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4644 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4645 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4646 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4647 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4648 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4649 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4650 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4651 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4652 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4653 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4654 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4655 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4656 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4657 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4658 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4659 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4660 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4661 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4662 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4663 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4664 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4665 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4666 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4667 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4668 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4669 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4670 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4671 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4672 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4673 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4674 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4675 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4676 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4677 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4678 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4679 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4680 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4681 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4682 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4683 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4684 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4685 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4686 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4687 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4688 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4689 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4690 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4691 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4692 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4693 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4694 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4695 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4696 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4697 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4698 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4699 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4700 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4701 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4702 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4703 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4704 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4705 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4706 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4707 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4708 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4709 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4710 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4711 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4712 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4713 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4714 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4715 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4716 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4717 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4718 x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4719 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4720 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4721 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4722 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4723 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4724 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4725 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4726 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4727 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4728 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4729 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4730 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4731 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4732 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4733 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4734 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4735 9bitdac_layout_0/8bitdac_layout_1/x1_vref5 9bitdac_layout_0/8bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4736 9bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4737 9bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4738 9bitdac_layout_1/switch_layout_0/dinb d8 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4739 9bitdac_layout_1/switch_layout_0/dinb d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4740 9bitdac_layout_1/x1_out_v 9bitdac_layout_1/switch_layout_0/dd x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4741 x2_out_v 9bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/x1_out_v 9bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4742 9bitdac_layout_1/x2_out_v 9bitdac_layout_1/switch_layout_0/dd x2_out_v 9bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4743 x2_out_v 9bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4744 9bitdac_layout_1/x1_vref5 9bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4745 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4746 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4747 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb d7 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4748 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4749 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4750 9bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4751 9bitdac_layout_1/8bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4752 9bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4753 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4754 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4755 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4756 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4757 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4758 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4759 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4760 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4761 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4762 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4763 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4764 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4765 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4766 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4767 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4768 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4769 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4770 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4771 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4772 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4773 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4774 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4775 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4776 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4777 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4778 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4779 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4780 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4781 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4782 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4783 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4784 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4785 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4786 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4787 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4788 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4789 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4790 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4791 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4792 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4793 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4794 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4795 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4796 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4797 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4798 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4799 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4800 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4801 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4802 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4803 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4804 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4805 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4806 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4807 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4808 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4809 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4810 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4811 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4812 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4813 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4814 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4815 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4816 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4817 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4818 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4819 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4820 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4821 x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4822 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4823 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4824 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4825 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4826 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4827 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4828 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4829 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4830 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4831 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4832 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4833 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4834 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4835 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4836 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4837 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4838 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4839 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4840 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4841 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4842 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4843 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4844 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4845 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4846 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4847 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4848 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4849 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4850 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4851 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4852 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4853 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4854 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4855 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4856 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4857 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4858 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4859 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4860 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4861 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4862 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4863 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4864 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4865 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4866 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4867 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4868 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4869 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4870 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4871 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4872 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4873 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4874 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4875 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4876 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4877 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4878 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4879 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4880 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4881 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4882 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4883 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4884 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4885 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4886 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4887 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4888 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4889 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4890 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4891 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4892 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4893 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4894 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4895 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4896 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4897 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4898 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4899 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4900 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4901 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4902 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4903 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4904 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4905 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4906 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4907 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4908 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4909 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4910 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4911 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4912 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4913 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4914 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4915 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4916 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4917 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4918 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4919 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4920 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4921 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4922 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4923 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4924 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4925 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4926 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4927 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4928 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4929 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4930 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4931 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4932 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4933 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4934 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4935 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4936 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4937 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4938 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4939 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4940 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4941 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4942 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4943 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4944 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4945 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4946 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4947 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4948 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4949 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4950 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4951 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4952 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4953 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4954 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4955 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4956 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4957 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4958 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4959 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4960 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4961 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4962 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4963 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4964 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4965 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4966 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4967 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4968 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4969 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4970 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4971 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4972 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4973 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4974 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4975 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4976 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4977 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4978 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4979 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4980 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4981 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4982 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4983 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4984 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4985 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4986 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4987 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4988 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X4989 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4990 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X4991 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4992 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4993 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X4994 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4995 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4996 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X4997 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X4998 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X4999 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5000 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5001 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5002 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5003 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5004 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5005 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5006 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5007 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5008 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5009 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5010 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5011 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5012 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5013 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5014 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5015 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5016 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5017 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5018 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5019 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5020 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5021 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5022 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5023 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5024 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5025 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5026 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5027 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5028 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5029 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5030 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5031 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5032 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5033 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5034 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5035 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5036 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5037 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5038 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5039 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5040 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5041 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5042 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5043 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5044 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5045 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5046 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5047 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5048 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5049 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5050 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5051 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5052 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5053 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5054 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5055 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5056 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5057 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5058 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5059 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5060 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5061 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5062 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5063 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5064 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5065 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5066 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5067 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5068 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5069 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5070 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5071 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5072 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5073 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5074 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5075 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5076 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5077 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5078 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5079 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5080 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5081 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5082 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5083 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5084 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5085 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5086 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5087 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5088 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5089 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5090 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5091 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5092 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5093 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5094 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5095 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5096 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5097 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5098 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5099 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5100 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5101 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5102 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5103 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5104 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5105 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5106 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5107 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5108 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5109 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5110 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5111 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5112 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5113 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5114 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5115 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5116 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5117 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5118 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5119 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5120 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5121 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5122 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5123 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5124 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5125 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5126 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5127 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5128 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5129 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5130 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5131 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5132 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5133 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5134 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5135 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5136 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5137 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5138 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5139 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5140 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5141 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5142 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5143 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5144 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5145 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5146 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5147 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5148 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5149 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5150 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5151 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5152 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5153 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5154 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5155 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5156 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5157 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5158 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5159 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5160 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5161 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5162 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5163 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5164 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5165 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5166 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5167 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5168 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5169 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5170 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5171 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5172 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5173 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5174 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5175 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5176 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5177 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5178 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5179 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5180 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5181 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5182 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5183 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5184 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5185 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5186 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5187 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5188 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5189 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5190 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5191 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5192 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5193 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5194 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5195 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5196 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5197 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5198 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5199 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5200 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5201 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5202 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5203 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5204 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5205 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5206 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5207 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5208 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5209 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5210 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5211 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5212 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5213 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5214 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5215 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5216 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5217 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5218 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5219 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5220 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5221 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5222 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5223 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5224 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5225 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5226 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5227 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5228 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5229 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5230 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5231 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5232 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5233 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5234 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5235 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5236 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5237 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5238 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5239 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5240 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5241 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5242 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5243 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5244 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5245 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5246 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5247 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5248 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5249 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5250 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5251 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5252 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5253 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5254 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5255 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5256 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5257 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5258 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5259 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5260 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5261 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5262 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5263 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5264 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5265 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5266 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5267 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5268 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5269 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5270 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5271 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5272 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5273 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5274 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5275 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5276 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5277 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5278 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5279 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5280 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5281 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5282 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5283 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5284 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5285 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5286 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5287 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5288 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5289 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5290 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5291 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5292 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5293 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5294 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5295 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5296 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5297 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5298 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5299 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5300 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5301 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5302 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5303 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5304 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5305 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5306 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5307 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5308 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5309 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5310 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5311 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5312 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5313 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5314 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5315 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5316 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5317 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5318 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5319 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5320 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5321 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5322 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5323 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5324 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5325 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5326 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5327 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5328 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5329 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5330 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5331 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5332 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5333 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5334 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5335 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5336 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5337 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5338 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5339 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5340 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5341 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5342 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5343 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5344 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5345 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5346 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5347 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5348 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5349 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5350 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5351 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5352 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5353 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5354 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5355 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5356 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5357 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5358 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5359 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5360 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5361 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5362 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5363 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5364 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5365 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5366 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5367 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5368 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5369 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5370 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5371 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5372 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5373 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5374 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5375 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5376 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5377 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5378 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5379 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5380 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5381 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5382 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5383 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5384 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5385 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5386 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5387 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5388 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5389 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5390 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5391 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5392 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5393 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5394 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5395 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5396 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5397 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5398 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5399 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5400 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5401 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5402 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5403 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5404 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5405 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5406 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5407 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5408 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5409 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5410 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5411 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5412 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5413 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5414 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5415 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5416 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5417 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5418 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5419 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5420 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5421 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5422 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5423 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5424 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5425 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5426 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5427 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5428 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5429 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5430 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5431 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5432 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5433 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5434 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5435 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5436 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5437 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5438 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5439 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5440 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5441 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5442 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5443 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5444 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5445 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5446 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5447 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5448 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5449 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5450 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5451 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5452 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5453 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5454 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5455 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5456 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5457 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5458 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5459 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5460 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5461 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5462 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5463 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5464 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5465 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5466 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5467 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5468 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5469 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5470 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5471 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5472 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5473 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5474 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5475 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5476 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5477 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5478 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5479 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5480 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5481 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5482 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5483 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5484 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5485 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5486 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5487 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5488 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5489 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5490 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5491 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5492 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5493 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5494 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5495 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5496 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5497 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5498 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5499 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5500 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5501 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5502 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5503 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5504 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5505 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5506 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5507 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5508 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5509 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5510 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5511 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5512 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5513 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5514 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5515 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5516 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5517 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5518 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5519 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5520 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5521 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5522 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5523 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5524 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5525 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5526 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5527 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5528 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5529 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5530 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5531 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5532 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5533 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5534 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5535 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5536 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5537 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5538 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5539 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5540 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5541 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5542 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5543 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5544 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5545 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5546 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5547 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5548 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5549 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5550 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5551 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5552 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5553 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5554 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5555 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5556 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5557 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5558 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5559 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5560 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5561 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5562 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5563 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5564 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5565 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5566 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5567 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5568 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5569 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5570 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5571 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5572 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5573 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5574 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5575 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5576 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5577 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5578 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5579 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5580 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5581 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5582 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5583 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5584 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5585 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5586 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5587 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5588 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5589 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5590 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5591 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5592 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5593 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5594 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5595 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5596 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5597 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5598 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5599 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5600 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5601 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5602 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5603 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5604 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5605 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5606 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5607 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5608 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5609 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5610 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5611 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5612 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5613 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5614 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5615 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5616 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5617 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5618 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5619 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5620 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5621 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5622 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5623 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5624 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5625 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5626 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5627 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5628 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5629 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5630 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5631 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5632 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5633 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5634 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5635 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5636 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5637 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5638 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5639 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5640 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5641 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5642 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5643 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5644 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5645 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5646 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5647 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5648 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5649 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5650 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5651 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5652 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5653 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5654 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5655 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5656 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5657 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5658 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5659 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5660 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5661 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5662 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5663 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5664 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5665 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5666 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5667 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5668 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5669 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5670 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5671 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5672 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5673 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5674 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5675 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5676 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5677 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5678 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5679 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5680 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5681 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5682 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5683 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5684 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5685 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5686 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5687 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5688 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5689 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5690 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5691 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5692 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5693 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5694 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5695 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5696 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5697 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5698 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5699 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5700 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5701 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5702 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5703 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5704 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5705 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5706 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5707 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5708 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5709 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5710 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5711 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5712 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5713 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5714 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5715 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5716 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5717 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5718 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5719 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5720 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5721 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5722 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5723 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5724 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5725 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5726 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5727 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5728 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5729 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5730 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5731 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5732 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5733 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5734 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5735 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5736 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5737 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5738 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5739 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5740 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5741 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5742 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5743 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5744 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5745 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5746 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5747 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5748 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5749 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5750 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5751 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5752 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5753 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5754 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5755 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5756 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5757 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5758 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5759 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5760 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5761 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5762 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5763 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5764 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5765 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5766 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5767 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5768 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5769 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5770 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5771 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5772 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5773 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5774 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5775 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5776 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5777 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5778 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5779 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5780 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5781 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5782 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5783 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5784 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5785 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5786 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5787 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5788 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5789 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5790 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5791 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5792 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5793 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5794 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5795 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5796 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5797 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5798 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5799 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5800 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5801 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5802 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5803 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5804 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5805 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5806 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5807 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5808 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5809 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5810 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5811 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5812 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5813 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5814 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5815 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5816 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5817 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5818 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5819 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5820 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5821 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5822 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5823 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5824 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5825 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5826 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5827 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5828 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5829 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5830 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5831 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5832 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5833 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5834 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5835 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5836 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5837 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5838 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5839 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5840 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5841 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5842 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5843 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5844 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5845 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5846 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5847 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5848 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5849 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5850 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5851 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5852 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5853 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5854 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5855 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5856 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5857 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5858 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5859 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5860 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5861 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5862 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5863 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5864 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5865 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5866 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5867 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5868 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5869 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5870 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5871 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5872 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5873 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5874 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5875 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5876 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5877 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5878 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5879 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5880 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5881 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5882 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5883 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5884 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5885 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5886 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5887 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5888 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5889 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5890 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5891 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5892 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5893 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5894 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5895 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5896 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5897 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5898 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5899 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5900 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5901 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5902 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5903 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5904 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5905 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5906 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5907 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5908 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5909 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5910 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5911 9bitdac_layout_1/8bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5912 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5913 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5914 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5915 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5916 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5917 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5918 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5919 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5920 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5921 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5922 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5923 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5924 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5925 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5926 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5927 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5928 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5929 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5930 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5931 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5932 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5933 9bitdac_layout_1/8bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5934 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5935 9bitdac_layout_1/8bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5936 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5937 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5938 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5939 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5940 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5941 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5942 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5943 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5944 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5945 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5946 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5947 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5948 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5949 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5950 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5951 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5952 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5953 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5954 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5955 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5956 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5957 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5958 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5959 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5960 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5961 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5962 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5963 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5964 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5965 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5966 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5967 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5968 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5969 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5970 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5971 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5972 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5973 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5974 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5975 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5976 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5977 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5978 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5979 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5980 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5981 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5982 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5983 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5984 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5985 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5986 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5987 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5988 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5989 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5990 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5991 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X5992 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X5993 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X5994 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5995 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5996 9bitdac_layout_1/8bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X5997 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X5998 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X5999 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6000 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6001 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6002 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6003 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6004 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6005 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6006 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6007 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6008 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6009 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6010 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6011 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6012 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6013 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6014 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6015 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6016 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6017 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6018 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6019 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6020 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6021 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6022 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6023 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6024 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6025 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6026 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6027 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6028 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6029 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6030 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6031 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6032 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6033 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6034 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6035 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6036 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6037 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6038 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6039 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6040 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6041 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6042 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6043 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6044 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6045 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6046 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6047 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6048 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6049 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6050 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6051 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6052 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6053 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6054 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6055 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6056 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6057 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6058 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6059 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6060 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6061 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6062 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6063 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6064 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6065 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6066 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6067 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6068 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6069 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6070 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6071 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6072 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6073 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6074 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6075 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6076 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6077 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6078 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6079 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6080 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6081 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6082 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6083 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6084 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6085 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6086 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6087 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6088 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6089 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6090 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6091 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6092 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6093 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6094 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6095 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6096 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6097 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6098 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6099 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6100 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6101 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6102 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6103 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6104 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6105 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6106 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6107 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6108 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6109 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6110 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6111 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6112 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6113 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6114 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6115 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6116 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6117 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6118 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6119 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6120 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6121 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6122 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6123 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6124 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6125 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6126 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6127 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6128 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6129 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6130 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6131 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6132 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6133 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6134 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6135 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6136 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6137 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6138 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6139 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6140 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6141 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6142 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6143 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6144 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6145 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6146 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6147 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6148 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6149 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6150 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6151 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6152 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6153 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6154 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6155 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6156 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6157 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6158 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6159 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6160 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6161 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6162 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6163 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6164 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6165 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6166 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6167 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6168 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6169 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6170 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6171 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6172 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6173 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6174 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6175 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6176 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6177 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6178 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6179 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6180 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6181 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6182 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6183 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6184 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6185 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6186 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6187 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6188 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6189 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6190 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6191 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6192 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6193 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6194 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6195 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6196 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6197 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6198 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6199 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6200 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6201 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6202 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6203 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6204 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6205 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6206 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6207 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6208 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6209 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6210 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6211 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6212 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6213 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6214 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6215 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6216 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6217 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6218 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6219 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6220 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6221 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6222 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6223 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6224 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6225 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6226 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6227 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6228 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6229 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6230 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6231 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6232 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6233 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6234 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6235 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6236 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6237 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6238 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6239 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6240 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6241 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6242 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6243 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6244 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6245 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6246 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6247 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6248 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6249 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6250 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6251 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6252 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6253 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6254 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6255 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6256 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6257 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6258 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6259 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6260 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6261 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6262 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6263 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6264 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6265 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6266 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6267 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6268 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6269 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6270 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6271 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6272 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6273 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6274 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6275 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6276 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6277 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6278 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6279 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6280 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6281 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6282 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6283 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6284 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6285 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6286 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6287 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6288 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6289 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6290 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6291 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6292 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6293 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6294 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6295 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6296 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6297 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6298 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6299 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6300 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6301 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6302 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6303 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6304 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6305 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6306 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6307 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6308 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6309 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6310 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6311 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6312 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6313 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6314 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6315 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6316 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6317 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6318 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6319 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6320 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6321 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6322 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6323 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6324 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6325 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6326 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6327 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6328 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6329 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6330 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6331 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6332 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6333 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6334 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6335 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6336 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6337 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6338 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6339 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6340 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6341 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6342 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6343 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6344 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6345 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6346 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6347 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6348 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6349 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6350 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6351 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6352 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6353 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6354 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6355 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6356 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6357 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6358 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6359 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6360 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6361 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6362 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6363 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6364 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6365 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6366 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6367 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6368 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6369 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6370 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6371 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6372 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6373 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6374 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6375 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6376 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6377 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6378 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6379 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6380 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6381 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6382 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6383 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6384 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6385 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6386 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6387 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6388 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6389 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6390 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6391 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6392 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6393 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6394 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6395 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6396 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6397 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6398 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6399 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6400 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6401 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6402 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6403 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6404 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6405 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6406 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6407 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6408 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6409 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6410 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6411 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6412 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6413 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6414 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6415 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6416 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6417 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6418 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6419 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6420 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6421 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6422 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6423 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6424 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6425 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6426 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6427 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6428 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6429 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6430 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6431 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6432 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6433 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6434 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6435 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6436 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6437 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6438 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6439 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6440 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6441 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6442 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6443 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6444 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6445 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6446 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6447 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6448 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6449 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6450 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6451 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6452 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6453 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6454 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6455 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6456 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6457 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6458 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6459 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6460 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6461 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6462 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6463 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6464 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6465 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6466 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6467 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6468 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6469 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6470 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6471 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6472 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6473 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6474 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6475 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6476 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6477 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6478 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6479 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6480 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6481 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6482 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6483 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6484 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6485 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6486 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6487 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6488 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6489 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6490 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6491 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6492 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6493 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6494 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6495 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6496 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6497 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6498 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6499 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6500 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6501 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6502 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6503 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6504 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6505 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6506 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6507 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6508 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6509 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6510 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6511 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6512 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6513 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6514 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6515 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6516 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6517 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6518 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6519 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6520 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6521 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6522 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6523 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6524 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6525 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6526 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6527 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6528 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6529 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6530 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6531 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6532 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6533 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6534 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6535 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6536 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6537 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6538 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6539 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6540 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6541 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6542 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6543 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6544 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6545 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6546 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6547 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6548 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6549 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6550 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6551 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6552 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6553 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6554 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6555 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6556 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6557 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6558 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6559 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6560 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6561 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6562 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6563 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6564 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6565 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6566 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6567 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6568 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6569 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6570 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6571 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6572 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6573 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6574 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6575 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6576 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6577 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6578 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6579 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6580 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6581 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6582 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6583 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6584 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6585 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6586 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6587 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6588 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6589 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6590 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6591 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6592 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6593 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6594 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6595 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6596 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6597 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6598 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6599 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6600 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6601 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6602 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6603 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6604 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6605 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6606 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6607 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6608 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6609 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6610 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6611 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6612 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6613 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6614 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6615 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6616 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6617 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6618 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6619 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6620 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6621 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6622 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6623 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6624 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6625 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6626 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6627 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6628 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6629 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6630 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6631 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6632 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6633 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6634 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6635 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6636 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6637 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6638 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6639 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6640 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6641 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6642 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6643 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6644 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6645 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6646 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6647 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6648 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6649 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6650 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6651 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6652 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6653 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6654 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6655 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6656 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6657 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6658 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6659 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6660 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6661 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6662 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6663 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6664 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6665 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6666 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6667 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6668 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6669 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6670 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6671 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6672 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6673 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6674 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6675 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6676 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6677 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6678 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6679 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6680 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6681 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6682 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6683 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6684 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6685 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6686 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6687 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6688 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6689 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6690 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6691 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6692 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6693 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6694 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6695 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6696 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6697 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6698 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6699 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6700 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6701 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6702 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6703 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6704 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6705 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6706 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6707 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6708 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6709 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6710 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6711 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6712 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6713 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6714 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6715 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6716 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6717 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6718 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6719 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6720 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6721 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6722 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6723 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6724 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6725 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6726 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6727 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6728 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6729 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6730 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6731 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6732 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6733 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6734 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6735 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6736 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6737 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6738 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6739 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6740 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6741 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6742 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6743 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6744 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6745 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6746 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6747 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6748 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6749 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6750 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6751 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6752 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6753 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6754 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6755 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6756 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6757 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6758 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6759 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6760 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6761 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6762 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6763 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6764 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6765 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6766 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6767 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6768 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6769 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6770 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6771 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6772 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6773 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6774 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6775 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6776 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6777 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6778 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6779 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6780 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6781 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6782 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6783 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6784 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6785 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6786 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6787 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6788 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6789 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6790 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6791 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6792 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6793 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6794 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6795 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6796 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6797 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6798 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6799 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6800 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6801 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6802 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6803 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6804 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6805 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6806 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6807 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6808 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6809 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6810 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6811 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6812 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6813 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6814 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6815 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6816 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6817 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6818 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6819 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6820 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6821 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6822 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6823 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6824 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6825 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6826 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6827 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6828 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6829 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6830 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6831 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6832 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6833 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6834 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6835 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6836 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6837 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6838 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6839 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6840 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6841 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6842 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6843 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6844 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6845 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6846 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6847 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6848 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6849 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6850 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6851 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6852 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6853 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6854 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6855 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6856 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6857 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6858 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6859 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6860 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6861 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6862 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6863 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6864 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6865 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6866 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6867 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6868 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6869 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6870 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6871 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6872 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6873 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6874 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6875 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6876 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6877 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6878 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6879 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6880 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6881 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6882 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6883 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6884 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6885 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6886 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6887 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6888 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6889 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6890 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6891 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6892 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6893 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6894 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6895 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6896 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6897 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6898 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6899 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6900 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6901 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6902 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6903 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6904 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6905 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6906 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6907 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6908 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6909 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6910 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6911 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6912 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6913 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6914 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6915 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6916 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6917 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6918 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6919 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6920 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6921 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6922 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6923 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6924 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6925 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6926 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6927 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6928 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6929 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6930 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6931 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6932 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6933 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6934 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6935 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6936 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6937 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6938 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6939 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6940 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6941 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6942 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6943 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6944 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6945 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6946 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6947 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6948 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6949 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6950 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6951 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6952 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6953 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6954 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6955 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6956 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6957 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6958 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6959 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X6960 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6961 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6962 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X6963 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6964 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6965 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6966 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6967 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6968 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6969 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6970 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6971 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6972 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6973 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6974 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6975 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6976 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6977 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6978 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6979 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6980 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6981 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6982 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6983 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6984 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6985 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6986 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6987 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6988 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6989 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6990 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6991 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6992 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X6993 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6994 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X6995 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6996 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6997 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X6998 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X6999 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7000 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7001 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7002 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7003 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7004 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7005 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7006 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7007 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7008 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7009 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7010 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7011 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7012 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7013 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7014 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7015 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7016 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7017 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7018 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7019 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7020 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7021 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7022 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7023 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7024 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7025 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7026 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7027 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7028 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7029 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7030 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7031 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7032 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7033 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7034 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7035 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7036 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7037 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7038 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7039 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7040 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7041 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7042 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7043 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7044 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7045 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7046 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7047 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7048 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7049 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7050 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7051 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7052 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7053 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7054 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7055 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7056 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7057 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7058 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7059 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7060 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7061 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7062 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7063 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7064 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7065 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7066 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7067 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7068 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7069 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7070 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7071 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7072 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7073 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7074 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7075 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7076 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7077 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7078 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7079 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7080 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7081 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7082 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7083 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7084 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7085 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7086 9bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7087 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7088 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7089 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7090 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7091 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7092 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7093 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7094 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7095 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7096 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7097 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7098 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7099 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7100 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7101 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7102 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7103 9bitdac_layout_1/8bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7104 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7105 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7106 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb d7 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7107 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7108 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7109 9bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7110 9bitdac_layout_1/8bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7111 9bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7112 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7113 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7114 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7115 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7116 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7117 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7118 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7119 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7120 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7121 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7122 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7123 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7124 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7125 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7126 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7127 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7128 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7129 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7130 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7131 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7132 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7133 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7134 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7135 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7136 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7137 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7138 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7139 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7140 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7141 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7142 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7143 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7144 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7145 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7146 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7147 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7148 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7149 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7150 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7151 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7152 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7153 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7154 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7155 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7156 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7157 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7158 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7159 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7160 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7161 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7162 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7163 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7164 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7165 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7166 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7167 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7168 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7169 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7170 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7171 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7172 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7173 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7174 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7175 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7176 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7177 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7178 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7179 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7180 9bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7181 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7182 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7183 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7184 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7185 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7186 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7187 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7188 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7189 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7190 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7191 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7192 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7193 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7194 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7195 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7196 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7197 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7198 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7199 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7200 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7201 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7202 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7203 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7204 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7205 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7206 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7207 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7208 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7209 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7210 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7211 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7212 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7213 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7214 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7215 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7216 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7217 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7218 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7219 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7220 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7221 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7222 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7223 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7224 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7225 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7226 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7227 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7228 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7229 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7230 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7231 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7232 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7233 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7234 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7235 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7236 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7237 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7238 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7239 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7240 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7241 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7242 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7243 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7244 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7245 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7246 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7247 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7248 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7249 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7250 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7251 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7252 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7253 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7254 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7255 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7256 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7257 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7258 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7259 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7260 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7261 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7262 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7263 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7264 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7265 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7266 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7267 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7268 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7269 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7270 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7271 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7272 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7273 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7274 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7275 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7276 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7277 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7278 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7279 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7280 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7281 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7282 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7283 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7284 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7285 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7286 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7287 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7288 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7289 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7290 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7291 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7292 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7293 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7294 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7295 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7296 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7297 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7298 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7299 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7300 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7301 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7302 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7303 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7304 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7305 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7306 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7307 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7308 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7309 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7310 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7311 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7312 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7313 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7314 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7315 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7316 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7317 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7318 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7319 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7320 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7321 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7322 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7323 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7324 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7325 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7326 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7327 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7328 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7329 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7330 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7331 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7332 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7333 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7334 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7335 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7336 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7337 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7338 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7339 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7340 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7341 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7342 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7343 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7344 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7345 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7346 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7347 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7348 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7349 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7350 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7351 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7352 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7353 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7354 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7355 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7356 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7357 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7358 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7359 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7360 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7361 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7362 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7363 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7364 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7365 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7366 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7367 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7368 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7369 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7370 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7371 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7372 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7373 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7374 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7375 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7376 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7377 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7378 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7379 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7380 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7381 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7382 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7383 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7384 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7385 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7386 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7387 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7388 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7389 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7390 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7391 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7392 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7393 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7394 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7395 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7396 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7397 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7398 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7399 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7400 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7401 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7402 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7403 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7404 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7405 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7406 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7407 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7408 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7409 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7410 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7411 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7412 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7413 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7414 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7415 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7416 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7417 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7418 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7419 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7420 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7421 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7422 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7423 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7424 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7425 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7426 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7427 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7428 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7429 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7430 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7431 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7432 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7433 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7434 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7435 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7436 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7437 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7438 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7439 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7440 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7441 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7442 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7443 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7444 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7445 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7446 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7447 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7448 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7449 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7450 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7451 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7452 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7453 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7454 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7455 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7456 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7457 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7458 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7459 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7460 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7461 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7462 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7463 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7464 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7465 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7466 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7467 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7468 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7469 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7470 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7471 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7472 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7473 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7474 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7475 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7476 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7477 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7478 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7479 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7480 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7481 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7482 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7483 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7484 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7485 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7486 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7487 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7488 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7489 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7490 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7491 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7492 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7493 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7494 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7495 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7496 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7497 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7498 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7499 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7500 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7501 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7502 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7503 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7504 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7505 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7506 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7507 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7508 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7509 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7510 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7511 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7512 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7513 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7514 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7515 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7516 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7517 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7518 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7519 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7520 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7521 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7522 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7523 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7524 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7525 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7526 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7527 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7528 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7529 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7530 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7531 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7532 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7533 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7534 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7535 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7536 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7537 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7538 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7539 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7540 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7541 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7542 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7543 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7544 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7545 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7546 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7547 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7548 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7549 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7550 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7551 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7552 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7553 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7554 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7555 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7556 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7557 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7558 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7559 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7560 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7561 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7562 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7563 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7564 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7565 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7566 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7567 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7568 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7569 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7570 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7571 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7572 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7573 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7574 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7575 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7576 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7577 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7578 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7579 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7580 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7581 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7582 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7583 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7584 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7585 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7586 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7587 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7588 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7589 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7590 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7591 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7592 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7593 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7594 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7595 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7596 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7597 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7598 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7599 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7600 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7601 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7602 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7603 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7604 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7605 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7606 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7607 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7608 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7609 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7610 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7611 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7612 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7613 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7614 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7615 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7616 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7617 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7618 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7619 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7620 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7621 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7622 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7623 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7624 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7625 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7626 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7627 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7628 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7629 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7630 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7631 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7632 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7633 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7634 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7635 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7636 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7637 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7638 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7639 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7640 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7641 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7642 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7643 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7644 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7645 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7646 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7647 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7648 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7649 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7650 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7651 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7652 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7653 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7654 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7655 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7656 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7657 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7658 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7659 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7660 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7661 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7662 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7663 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7664 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7665 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7666 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7667 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7668 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7669 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7670 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7671 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7672 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7673 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7674 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7675 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7676 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7677 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7678 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7679 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7680 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7681 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7682 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7683 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7684 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7685 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7686 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7687 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7688 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7689 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7690 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7691 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7692 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7693 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7694 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7695 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7696 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7697 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7698 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7699 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7700 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7701 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7702 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7703 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7704 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7705 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7706 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7707 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7708 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7709 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7710 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7711 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7712 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7713 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7714 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7715 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7716 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7717 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7718 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7719 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7720 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7721 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7722 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7723 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7724 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7725 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7726 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7727 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7728 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7729 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7730 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7731 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7732 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7733 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7734 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7735 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7736 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7737 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7738 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7739 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7740 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7741 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7742 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7743 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7744 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7745 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7746 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7747 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7748 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7749 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7750 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7751 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7752 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7753 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7754 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7755 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7756 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7757 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7758 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7759 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7760 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7761 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7762 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7763 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7764 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7765 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7766 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7767 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7768 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7769 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7770 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7771 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7772 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7773 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7774 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7775 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7776 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7777 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7778 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7779 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7780 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7781 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7782 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7783 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7784 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7785 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7786 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7787 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7788 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7789 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7790 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7791 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7792 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7793 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7794 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7795 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7796 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7797 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7798 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7799 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7800 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7801 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7802 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7803 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7804 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7805 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7806 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7807 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7808 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7809 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7810 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7811 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7812 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7813 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7814 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7815 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7816 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7817 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7818 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7819 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7820 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7821 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7822 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7823 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7824 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7825 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7826 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7827 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7828 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7829 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7830 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7831 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7832 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7833 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7834 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7835 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7836 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7837 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7838 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7839 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7840 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7841 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7842 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7843 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7844 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7845 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7846 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7847 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7848 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7849 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7850 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7851 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7852 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7853 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7854 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7855 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7856 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7857 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7858 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7859 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7860 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7861 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7862 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7863 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7864 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7865 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7866 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7867 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7868 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7869 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7870 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7871 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7872 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7873 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7874 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7875 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7876 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7877 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7878 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7879 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7880 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7881 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7882 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7883 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7884 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7885 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7886 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7887 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7888 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7889 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7890 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7891 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7892 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7893 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7894 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7895 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7896 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7897 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7898 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7899 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7900 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7901 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7902 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7903 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7904 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7905 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7906 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7907 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7908 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7909 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7910 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7911 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7912 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7913 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7914 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7915 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7916 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7917 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7918 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7919 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7920 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7921 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7922 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7923 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7924 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7925 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7926 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7927 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7928 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7929 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7930 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7931 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7932 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7933 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7934 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7935 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7936 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7937 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7938 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7939 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7940 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7941 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7942 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7943 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7944 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7945 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7946 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7947 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7948 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7949 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7950 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7951 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7952 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7953 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7954 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7955 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7956 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7957 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7958 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7959 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7960 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7961 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7962 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7963 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7964 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7965 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7966 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7967 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7968 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7969 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7970 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7971 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7972 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7973 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7974 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7975 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7976 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7977 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7978 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7979 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7980 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7981 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7982 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7983 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7984 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7985 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7986 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7987 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X7988 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7989 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7990 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X7991 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X7992 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X7993 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7994 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7995 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X7996 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7997 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7998 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X7999 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8000 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8001 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8002 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8003 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8004 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8005 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8006 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8007 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8008 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8009 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8010 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8011 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8012 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8013 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8014 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8015 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8016 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8017 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8018 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8019 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8020 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8021 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8022 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8023 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8024 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8025 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8026 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8027 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8028 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8029 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8030 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8031 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8032 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8033 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8034 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8035 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8036 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8037 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8038 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8039 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8040 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8041 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8042 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8043 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8044 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8045 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8046 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8047 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8048 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8049 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8050 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8051 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8052 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8053 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8054 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8055 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8056 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8057 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8058 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8059 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8060 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8061 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8062 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8063 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8064 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8065 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8066 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8067 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8068 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8069 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8070 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8071 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8072 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8073 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8074 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8075 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8076 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8077 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8078 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8079 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8080 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8081 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8082 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8083 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8084 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8085 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8086 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8087 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8088 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8089 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8090 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8091 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8092 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8093 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8094 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8095 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8096 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8097 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8098 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8099 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8100 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8101 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8102 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8103 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8104 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8105 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8106 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8107 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8108 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8109 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8110 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8111 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8112 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8113 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8114 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8115 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8116 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8117 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8118 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8119 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8120 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8121 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8122 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8123 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8124 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8125 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8126 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8127 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8128 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8129 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8130 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8131 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8132 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8133 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8134 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8135 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8136 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8137 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8138 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8139 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8140 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8141 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8142 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8143 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8144 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8145 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8146 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8147 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8148 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8149 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8150 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8151 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8152 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8153 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8154 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8155 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8156 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8157 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8158 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8159 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8160 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8161 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8162 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8163 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8164 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8165 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8166 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8167 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8168 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8169 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8170 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8171 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8172 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8173 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8174 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8175 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8176 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8177 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8178 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8179 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8180 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8181 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8182 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8183 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8184 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8185 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8186 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8187 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8188 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8189 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8190 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8191 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8192 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8193 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8194 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8195 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8196 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8197 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8198 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8199 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8200 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8201 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8202 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8203 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8204 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8205 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8206 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8207 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8208 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8209 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8210 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8211 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8212 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8213 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8214 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8215 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8216 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8217 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8218 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8219 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8220 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8221 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8222 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8223 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8224 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8225 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8226 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8227 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8228 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8229 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8230 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8231 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8232 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8233 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8234 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8235 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8236 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8237 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8238 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8239 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8240 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8241 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8242 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8243 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8244 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8245 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8246 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8247 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8248 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8249 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8250 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8251 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8252 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8253 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8254 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8255 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8256 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8257 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8258 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8259 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8260 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8261 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8262 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8263 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8264 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8265 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8266 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8267 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8268 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8269 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8270 9bitdac_layout_1/8bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8271 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8272 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8273 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8274 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8275 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8276 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8277 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8278 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8279 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8280 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8281 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8282 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8283 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8284 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8285 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8286 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8287 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8288 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8289 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb d6 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8290 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8291 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8292 9bitdac_layout_1/8bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8293 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8294 9bitdac_layout_1/8bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8295 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8296 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8297 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8298 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8299 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8300 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8301 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8302 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8303 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8304 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8305 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8306 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8307 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8308 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8309 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8310 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8311 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8312 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8313 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8314 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8315 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8316 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8317 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8318 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8319 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8320 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8321 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8322 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8323 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8324 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8325 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8326 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8327 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8328 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8329 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8330 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8331 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8332 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8333 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8334 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8335 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8336 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8337 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8338 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8339 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8340 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8341 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8342 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8343 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8344 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8345 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8346 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8347 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8348 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8349 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8350 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8351 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8352 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8353 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8354 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8355 9bitdac_layout_1/8bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8356 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8357 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8358 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8359 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8360 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8361 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8362 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8363 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8364 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8365 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8366 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8367 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8368 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8369 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8370 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8371 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8372 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8373 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8374 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8375 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8376 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8377 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8378 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8379 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8380 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8381 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8382 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8383 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8384 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8385 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8386 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8387 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8388 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8389 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8390 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8391 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8392 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8393 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8394 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8395 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8396 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8397 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8398 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8399 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8400 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8401 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8402 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8403 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8404 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8405 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8406 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8407 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8408 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8409 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8410 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8411 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8412 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8413 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8414 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8415 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8416 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8417 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8418 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8419 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8420 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8421 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8422 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8423 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8424 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8425 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8426 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8427 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8428 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8429 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8430 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8431 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8432 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8433 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8434 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8435 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8436 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8437 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8438 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8439 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8440 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8441 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8442 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8443 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8444 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8445 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8446 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8447 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8448 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8449 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8450 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8451 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8452 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8453 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8454 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8455 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8456 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8457 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8458 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8459 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8460 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8461 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8462 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8463 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8464 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8465 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8466 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8467 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8468 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8469 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8470 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8471 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8472 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8473 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8474 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8475 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8476 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8477 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8478 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8479 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8480 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8481 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8482 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8483 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8484 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8485 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8486 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8487 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8488 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8489 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8490 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8491 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8492 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8493 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8494 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8495 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8496 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8497 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8498 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8499 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8500 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8501 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8502 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8503 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8504 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8505 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8506 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8507 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8508 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8509 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8510 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8511 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8512 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8513 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8514 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8515 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8516 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8517 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8518 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8519 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8520 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8521 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8522 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8523 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8524 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8525 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8526 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8527 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8528 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8529 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8530 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8531 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8532 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8533 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8534 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8535 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8536 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8537 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8538 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8539 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8540 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8541 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8542 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8543 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8544 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8545 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8546 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8547 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8548 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8549 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8550 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8551 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8552 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8553 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8554 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8555 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8556 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8557 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8558 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8559 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8560 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8561 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8562 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8563 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8564 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8565 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8566 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8567 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8568 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8569 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8570 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8571 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8572 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8573 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8574 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8575 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8576 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8577 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8578 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8579 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8580 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8581 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8582 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8583 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8584 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8585 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8586 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8587 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8588 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8589 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8590 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8591 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8592 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8593 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8594 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8595 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8596 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8597 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8598 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8599 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8600 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8601 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8602 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8603 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8604 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8605 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8606 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8607 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8608 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8609 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8610 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8611 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8612 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8613 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8614 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8615 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8616 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8617 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8618 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8619 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8620 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8621 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8622 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8623 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8624 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8625 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8626 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8627 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8628 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8629 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8630 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8631 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8632 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8633 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8634 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8635 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8636 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8637 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8638 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8639 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8640 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8641 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8642 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8643 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8644 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8645 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8646 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8647 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8648 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8649 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8650 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8651 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8652 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8653 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8654 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8655 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8656 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8657 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8658 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8659 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8660 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8661 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8662 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8663 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8664 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8665 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8666 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8667 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8668 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8669 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8670 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8671 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8672 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8673 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8674 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8675 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8676 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8677 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8678 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8679 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8680 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8681 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8682 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8683 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8684 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8685 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8686 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8687 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8688 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8689 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8690 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8691 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8692 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8693 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8694 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8695 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8696 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8697 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8698 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8699 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8700 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8701 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8702 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8703 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8704 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8705 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8706 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8707 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8708 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8709 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8710 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8711 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8712 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8713 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8714 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8715 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8716 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8717 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8718 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8719 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8720 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8721 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8722 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8723 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8724 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8725 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8726 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8727 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8728 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8729 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8730 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8731 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8732 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8733 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8734 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8735 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8736 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8737 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8738 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8739 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8740 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8741 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8742 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8743 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8744 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8745 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8746 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8747 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8748 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8749 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8750 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8751 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8752 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8753 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8754 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8755 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8756 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8757 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8758 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8759 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8760 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8761 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8762 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8763 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8764 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8765 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8766 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8767 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8768 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8769 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8770 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8771 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8772 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8773 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8774 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8775 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8776 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8777 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8778 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8779 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8780 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8781 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8782 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8783 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8784 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8785 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8786 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8787 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8788 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8789 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8790 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8791 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8792 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8793 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8794 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8795 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8796 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8797 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8798 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8799 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8800 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8801 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8802 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8803 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8804 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8805 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8806 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8807 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8808 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8809 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8810 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8811 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8812 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8813 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8814 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8815 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8816 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8817 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8818 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8819 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8820 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8821 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8822 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8823 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8824 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8825 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8826 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8827 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8828 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8829 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8830 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8831 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8832 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8833 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8834 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8835 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8836 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8837 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8838 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8839 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8840 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8841 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8842 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8843 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8844 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8845 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8846 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8847 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8848 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8849 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8850 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8851 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8852 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8853 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8854 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8855 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8856 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8857 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8858 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8859 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8860 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8861 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8862 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8863 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8864 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8865 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8866 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8867 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8868 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8869 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8870 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8871 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8872 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8873 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8874 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8875 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8876 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8877 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8878 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8879 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8880 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8881 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8882 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8883 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8884 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8885 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8886 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8887 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8888 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8889 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8890 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8891 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8892 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8893 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8894 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8895 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8896 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8897 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8898 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8899 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8900 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8901 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8902 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8903 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8904 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8905 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8906 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8907 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8908 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8909 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8910 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8911 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8912 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8913 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8914 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8915 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8916 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8917 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8918 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8919 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8920 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8921 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8922 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8923 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8924 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8925 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8926 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8927 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8928 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8929 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8930 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8931 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8932 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8933 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8934 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8935 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8936 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8937 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8938 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8939 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8940 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8941 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8942 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8943 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8944 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8945 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8946 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8947 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8948 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8949 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8950 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8951 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8952 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8953 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8954 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8955 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8956 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8957 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8958 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8959 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8960 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8961 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8962 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8963 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8964 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8965 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8966 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X8967 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8968 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X8969 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8970 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8971 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8972 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8973 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8974 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8975 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8976 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8977 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8978 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8979 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8980 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8981 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8982 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8983 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8984 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8985 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8986 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8987 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8988 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8989 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8990 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8991 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8992 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8993 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8994 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8995 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X8996 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X8997 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X8998 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X8999 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9000 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9001 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9002 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9003 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9004 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9005 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9006 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9007 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9008 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9009 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9010 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9011 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9012 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9013 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9014 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9015 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9016 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9017 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9018 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9019 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9020 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9021 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9022 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9023 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9024 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9025 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9026 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9027 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9028 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9029 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9030 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9031 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9032 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9033 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9034 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9035 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9036 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9037 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9038 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9039 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9040 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9041 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9042 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9043 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9044 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9045 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9046 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9047 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9048 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9049 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9050 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9051 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9052 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9053 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9054 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9055 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9056 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9057 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9058 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9059 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9060 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9061 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9062 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9063 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9064 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9065 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9066 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9067 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9068 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9069 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9070 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9071 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9072 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9073 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9074 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9075 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9076 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9077 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9078 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9079 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9080 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9081 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9082 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9083 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9084 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9085 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9086 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9087 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9088 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9089 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9090 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9091 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9092 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9093 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9094 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9095 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9096 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9097 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9098 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9099 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9100 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9101 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9102 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9103 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9104 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9105 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9106 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9107 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9108 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9109 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9110 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9111 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9112 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9113 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9114 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9115 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9116 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9117 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9118 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9119 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9120 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9121 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9122 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9123 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9124 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9125 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9126 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9127 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9128 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9129 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9130 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9131 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9132 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9133 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9134 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9135 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9136 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9137 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9138 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9139 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9140 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9141 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9142 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9143 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9144 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9145 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9146 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9147 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9148 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9149 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9150 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9151 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9152 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9153 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9154 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9155 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9156 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9157 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9158 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9159 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9160 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9161 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9162 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9163 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9164 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9165 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9166 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9167 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9168 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9169 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9170 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9171 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9172 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9173 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9174 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9175 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9176 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9177 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9178 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9179 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9180 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9181 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9182 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9183 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9184 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9185 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9186 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9187 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9188 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9189 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9190 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9191 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9192 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9193 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9194 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9195 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9196 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9197 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9198 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9199 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9200 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9201 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9202 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9203 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9204 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9205 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9206 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9207 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9208 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9209 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9210 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9211 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9212 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9213 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9214 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9215 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9216 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9217 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9218 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9219 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9220 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9221 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9222 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9223 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9224 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9225 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9226 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9227 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9228 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9229 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9230 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9231 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9232 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9233 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9234 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9235 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9236 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9237 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9238 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9239 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9240 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9241 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9242 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9243 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9244 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9245 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9246 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9247 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9248 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9249 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9250 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9251 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9252 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9253 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9254 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9255 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9256 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9257 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9258 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9259 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9260 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9261 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9262 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9263 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9264 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9265 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9266 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9267 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9268 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9269 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9270 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9271 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9272 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9273 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9274 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9275 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9276 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9277 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9278 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9279 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9280 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9281 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9282 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9283 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9284 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9285 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9286 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9287 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9288 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9289 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9290 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9291 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9292 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9293 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9294 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9295 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9296 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9297 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9298 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9299 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9300 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9301 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9302 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9303 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9304 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9305 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9306 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9307 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9308 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9309 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9310 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9311 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9312 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9313 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9314 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9315 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9316 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9317 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9318 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9319 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9320 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9321 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9322 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9323 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9324 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9325 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9326 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9327 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9328 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9329 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9330 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9331 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9332 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9333 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9334 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9335 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9336 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9337 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9338 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9339 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9340 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9341 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9342 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9343 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9344 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9345 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9346 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9347 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9348 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9349 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9350 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9351 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9352 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9353 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9354 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9355 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9356 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9357 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9358 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9359 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9360 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9361 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9362 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9363 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9364 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9365 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9366 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9367 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9368 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9369 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9370 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9371 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9372 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9373 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9374 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9375 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9376 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9377 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9378 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9379 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9380 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9381 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9382 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9383 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9384 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9385 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9386 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9387 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9388 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9389 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9390 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9391 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9392 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9393 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9394 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_0/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9395 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9396 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9397 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9398 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9399 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9400 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9401 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9402 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9403 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9404 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9405 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9406 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9407 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9408 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9409 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9410 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9411 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9412 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9413 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9414 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9415 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9416 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9417 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9418 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9419 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9420 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9421 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9422 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9423 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9424 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9425 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9426 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9427 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9428 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9429 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9430 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_0/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9431 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9432 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9433 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9434 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9435 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9436 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9437 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9438 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_0/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9439 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9440 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9441 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9442 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9443 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9444 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9445 inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9446 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_1/dinb inp2 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9447 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9448 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9449 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 0 0 sky130_fd_pr__nfet_01v8 w=0.61 l=0.15
X9450 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9451 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9452 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_583_327# sky130_fd_pr__pfet_01v8 w=1.21 l=0.15
X9453 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dd 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/w_908_86# sky130_fd_pr__pfet_01v8 w=1.20 l=0.15
X9454 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_out_v 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/switch_layout_2/dinb 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_vout 0 sky130_fd_pr__nfet_01v8 w=0.60 l=0.15
X9455 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9456 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp2 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9457 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x1_inp1 0 sky130_fd_pr__res_generic_nd w=0.27 l=1.24
X9458 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/2bitdac_layout_1/x2_inp1 inp2 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9459 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/3bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9460 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9461 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
X9462 9bitdac_layout_1/8bitdac_layout_1/x1_vref5 9bitdac_layout_1/8bitdac_layout_1/x2_vref1 0 sky130_fd_pr__res_generic_nd w=0.29 l=0.65
C0 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/x2_vref1 12.72fF
C1 9bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 19.77fF
C2 vdd d2 8.96fF
C3 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 2.44fF
C4 d6 d0 28.63fF
C5 d4 d2 20.08fF
C6 d5 d7 4.02fF
C7 vdd d1 42.81fF
C8 d2 d1 49.96fF
C9 d4 d1 7.44fF
C10 d2 d0 16.85fF
C11 vdd d3 6.90fF
C12 d2 d3 67.70fF
C13 d4 d3 129.84fF
C14 d1 d0 179.55fF
C15 d3 d0 6.80fF
C16 9bitdac_layout_1/x2_vref1 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 3.29fF
C17 9bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/x1_out_v 3.29fF
C18 9bitdac_layout_0/8bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 2.44fF
C19 x2_vref1 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 8.21fF
C20 d5 d2 3.34fF
C21 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/x2_vref1 12.72fF
C22 d5 d4 95.86fF
C23 x2_vref1 9bitdac_layout_1/x1_out_v 5.86fF
C24 d6 d1 15.27fF
C25 d5 d0 11.54fF
C26 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 9bitdac_layout_1/8bitdac_layout_0/x1_out_v 2.44fF
C27 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/x2_vref1 12.72fF
C28 d2 d1 49.96fF
C29 9bitdac_layout_0/8bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_out_v 12.72fF
C30 9bitdac_layout_1/8bitdac_layout_1/x2_vref1 9bitdac_layout_1/x1_out_v 3.09fF
C31 vdd d2 8.89fF
C32 d2 d3 67.70fF
C33 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 9bitdac_layout_1/x1_out_v 34.19fF
C34 d7 d6 23.66fF
C35 d4 d2 20.08fF
C36 d3 d1 36.27fF
C37 9bitdac_layout_0/x2_vref1 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_out_v 19.77fF
C38 vdd d0 53.48fF
C39 9bitdac_layout_0/8bitdac_layout_1/x1_out_v 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_out_v 2.44fF
C40 d5 d6 56.74fF
C41 d2 d0 16.90fF
C42 x2_vref1 9bitdac_layout_1/8bitdac_layout_1/x1_out_v 3.14fF
C43 d4 d0 5.09fF
C44 9bitdac_layout_0/8bitdac_layout_1/x2_vref1 9bitdac_layout_0/x1_out_v 3.09fF
C45 d5 d2 3.34fF
C46 d5 d1 5.05fF
C47 d5 d3 29.02fF
C48 9bitdac_layout_0/8bitdac_layout_1/x1_out_v 9bitdac_layout_0/x1_out_v 34.19fF
C49 d4 d6 22.94fF
C50 vdd 0 1922.01fF
C51 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C52 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C53 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C54 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C55 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 2.08fF
C56 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C57 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C58 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C59 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C60 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C61 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C62 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C63 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C64 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 2.08fF
C65 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C66 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C67 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C68 9bitdac_layout_1/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C69 9bitdac_layout_1/x1_vref5 0 2.19fF
C70 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C71 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C72 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C73 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C74 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 2.08fF
C75 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C76 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C77 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C78 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C79 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C80 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C81 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C82 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C83 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 2.08fF
C84 d0 0 858.43fF
C85 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C86 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C87 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C88 9bitdac_layout_1/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C89 d5 0 506.12fF
C90 d6 0 310.51fF
C91 d7 0 169.86fF
C92 x1_vref5 0 2.09fF
C93 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C94 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C95 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C96 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C97 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/x1_vref5 0 2.08fF
C98 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C99 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C100 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C101 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C102 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C103 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C104 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C105 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C106 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/x1_vref5 0 2.08fF
C107 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C108 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C109 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C110 9bitdac_layout_0/8bitdac_layout_1/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C111 9bitdac_layout_0/x1_vref5 0 2.19fF
C112 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C113 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C114 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C115 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C116 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/x1_vref5 0 2.08fF
C117 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C118 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C119 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C120 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_1/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C121 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C122 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C123 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C124 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_1/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF
C125 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/x1_vref5 0 2.08fF
C126 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_1/x1_vref5 0 2.13fF
C127 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_1/4bitdac_layout_0/x1_vref5 0 2.13fF
C128 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_1/x1_vref5 0 2.13fF
C129 9bitdac_layout_0/8bitdac_layout_0/7bitdac_layout_0/6bitdac_layout_0/5bitdac_layout_0/4bitdac_layout_0/x1_vref5 0 2.13fF


X9463 out_v 0 sky130_fd_pr__cap_mim_m3_1 W=25 L=25 MF=1

V1 vdd 0 dc 3.3V
V2 d0 0 PULSE 0 1.8 0ns 1p 1p 5u 10u
V3 d1 0 PULSE 0 1.8 0ns 1p 1p 10u 20u
V4 inp2 0 dc 0V
V5 inp1 0 dc 3.3V
V6 d2 0 PULSE 0 1.8 0ns 1p 1p 20u 40u
V7 d3 0 PULSE 0 1.8 0ns 1p 1p 40u 80u
V8 d4 0 PULSE 0 1.8 0ns 1p 1p 80u 160u
V9 d5 0 PULSE 0 1.8 0ns 1p 1p 160u 320u
V10 d6 0 PULSE 0 1.8 0 1p 1p 320u 640u
V11 d7 0 PULSE 0 1.8 0 1p 1p 640u 1280u
V12 d8 0 PULSE 0 1.8 0 1p 1p 1280u 2560u
V13 d9 0 PULSE 0 1.8 0 1p 1p 2560u 5120u

.tran 2u 5120u
.control
run 
plot d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 out_v
plot out_v
.endc
.end
