magic
tech sky130A
magscale 1 2
timestamp 1640022418
<< locali >>
rect 143604 52756 173468 52758
rect 143604 52718 198410 52756
rect 120322 52714 198410 52718
rect 120322 52674 143648 52714
rect 173454 52712 198410 52714
rect 97118 52582 97268 52584
rect 120322 52582 120364 52674
rect 97118 52576 120364 52582
rect 97118 52542 97135 52576
rect 97169 52542 120364 52576
rect 97118 52530 120364 52542
rect 97118 52528 120360 52530
rect 96280 52462 96342 52466
rect 98716 52462 98882 52466
rect 71454 52454 85650 52456
rect 94858 52454 96112 52456
rect 69398 52450 96112 52454
rect 67656 52446 67710 52448
rect 68402 52446 96112 52450
rect 67656 52434 96057 52446
rect 67656 52400 67662 52434
rect 67696 52412 96057 52434
rect 96091 52412 96112 52446
rect 96258 52452 98882 52462
rect 96258 52418 96285 52452
rect 96319 52418 98882 52452
rect 96258 52414 98882 52418
rect 96258 52412 97512 52414
rect 67696 52408 96112 52412
rect 67696 52406 71464 52408
rect 85622 52406 96112 52408
rect 67696 52402 69446 52406
rect 96040 52402 96108 52406
rect 96280 52404 96342 52412
rect 67696 52400 68450 52402
rect 67656 52398 68450 52400
rect 67656 52392 67710 52398
rect 97118 52322 97184 52334
rect 97118 52288 97135 52322
rect 97169 52288 97184 52322
rect 796 51892 854 51954
rect 67650 51664 67710 51674
rect 67650 51630 67664 51664
rect 67698 51630 67710 51664
rect 67650 51616 67710 51630
rect 67658 47534 67700 51616
rect 67658 41838 67702 47534
rect 67658 41806 67704 41838
rect 67660 36140 67704 41806
rect 67658 36110 67704 36140
rect 67658 24756 67702 36110
rect 97118 29332 97184 52288
rect 98820 52248 98878 52414
rect 98822 51746 98878 52248
rect 97112 28286 97184 29332
rect 198360 29304 198410 52712
rect 198360 29290 198412 29304
rect 198362 28628 198412 29290
rect 96494 28216 97184 28286
rect 198360 28592 198412 28628
rect 93744 28088 93994 28136
rect 93748 27571 93830 28088
rect 191874 28014 192000 28028
rect 191874 27918 192008 28014
rect 191876 27914 191984 27918
rect 93748 27537 93776 27571
rect 93810 27537 93830 27571
rect 93748 27504 93830 27537
rect 191880 27848 191942 27914
rect 191880 27404 191938 27848
rect 191880 27370 191891 27404
rect 191925 27370 191938 27404
rect 191880 27360 191938 27370
rect 194514 27280 194548 28140
rect 198360 27710 198410 28592
rect 198528 27444 198610 27446
rect 198526 27426 198772 27444
rect 198526 27392 198542 27426
rect 198576 27392 198772 27426
rect 198526 27380 198772 27392
rect 198528 27374 198610 27380
rect 93748 27185 93834 27210
rect 93748 27151 93774 27185
rect 93808 27151 93834 27185
rect 93748 26488 93834 27151
rect 192100 27050 192152 27056
rect 191880 27037 192152 27050
rect 191880 27003 191892 27037
rect 191926 27003 192152 27037
rect 194514 27012 194552 27280
rect 196098 27218 196190 27310
rect 191880 26992 192152 27003
rect 93752 26436 93830 26488
rect 93748 26284 93830 26436
rect 67658 24732 67704 24756
rect 67660 19046 67704 24732
rect 67658 16746 67704 19046
rect 67658 16720 67706 16746
rect 67660 14448 67706 16720
rect 67660 13050 67708 14448
rect 67658 13028 67708 13050
rect 67658 11654 67706 13028
rect 67658 11630 67708 11654
rect 67660 7450 67708 11630
rect 67658 7430 67708 7450
rect 67658 6042 67706 7430
rect 67656 6030 67706 6042
rect 67656 4634 67704 6030
rect 67654 4622 67704 4634
rect 67654 3230 67702 4622
rect 67862 3504 68030 3528
rect 67860 3490 68030 3504
rect 67860 3286 67908 3490
rect 67654 2942 67704 3230
rect 68032 2942 68084 3090
rect 67654 2894 68084 2942
rect 67654 2890 68082 2894
rect 93748 2452 93800 26284
rect 165990 3266 166048 3372
rect 93742 2428 93800 2452
rect 115660 2438 115708 2446
rect 68750 82 68816 100
rect 68750 48 68764 82
rect 68798 48 68816 82
rect 68750 30 68816 48
rect 68750 28 68818 30
rect 68760 18 68818 28
rect 68762 -226 68818 18
rect 68762 -1852 68808 -226
rect 68758 -1920 68808 -1852
rect 71804 -1830 71850 212
rect 75294 -1714 75370 414
rect 78572 -1620 78624 578
rect 81708 -1502 81778 784
rect 85106 -1290 85168 968
rect 90368 452 90440 1178
rect 90360 344 90440 452
rect 90360 -1042 90438 344
rect 93742 -868 93786 2428
rect 115660 2404 115667 2438
rect 115701 2404 115708 2438
rect 115660 2396 115708 2404
rect 112774 1876 112838 1984
rect 112776 1866 112838 1876
rect 112776 1832 112790 1866
rect 112824 1860 112838 1866
rect 112824 1832 112840 1860
rect 112776 1826 112840 1832
rect 112776 1824 112838 1826
rect 109158 1705 109194 1706
rect 109158 1671 109159 1705
rect 109193 1671 109194 1705
rect 109158 1670 109194 1671
rect 105668 1457 105754 1500
rect 105668 1423 105690 1457
rect 105724 1423 105754 1457
rect 105668 1396 105754 1423
rect 102398 1231 102442 1234
rect 102398 1197 102403 1231
rect 102437 1197 102442 1231
rect 192100 1198 192152 26992
rect 194506 26798 194556 27012
rect 194506 26794 195966 26798
rect 198380 26794 198430 26960
rect 194506 26740 198430 26794
rect 194506 26732 198422 26740
rect 195560 26728 198422 26732
rect 102398 1194 102442 1197
rect 99338 232 99406 1136
rect 102376 965 102454 1006
rect 102376 931 102403 965
rect 102437 931 102454 965
rect 105658 1001 105738 1032
rect 109150 1018 109200 1020
rect 105658 967 105680 1001
rect 105714 967 105738 1001
rect 105658 952 105738 967
rect 109148 1007 109200 1018
rect 109148 973 109157 1007
rect 109191 973 109200 1007
rect 109148 960 109200 973
rect 112780 968 112838 996
rect 102376 472 102454 931
rect 99338 -764 99402 232
rect 102376 -645 102444 472
rect 105670 134 105714 952
rect 102376 -679 102391 -645
rect 102425 -679 102444 -645
rect 102376 -714 102444 -679
rect 105672 -750 105714 134
rect 109148 -684 109196 960
rect 112780 934 112794 968
rect 112828 934 112838 968
rect 112780 228 112838 934
rect 141138 968 141176 970
rect 141138 934 141140 968
rect 141174 934 141176 968
rect 141138 932 141176 934
rect 115634 898 115734 928
rect 115634 864 115667 898
rect 115701 864 115734 898
rect 115634 458 115734 864
rect 112776 58 112838 228
rect 115628 274 115734 458
rect 112776 -660 112834 58
rect 99338 -798 99348 -764
rect 99382 -798 99402 -764
rect 99338 -808 99402 -798
rect 105670 -766 105740 -750
rect 105670 -800 105683 -766
rect 105717 -800 105740 -766
rect 109148 -760 109200 -684
rect 112776 -694 112792 -660
rect 112826 -694 112834 -660
rect 115628 -692 115728 274
rect 112776 -710 112834 -694
rect 115626 -724 115728 -692
rect 115626 -730 115669 -724
rect 109148 -794 109156 -760
rect 109190 -794 109200 -760
rect 115628 -758 115669 -730
rect 115703 -758 115728 -724
rect 115628 -776 115728 -758
rect 109148 -800 109200 -794
rect 105670 -814 105740 -800
rect 192090 -830 192162 1198
rect 192090 -860 192158 -830
rect 188778 -868 192158 -860
rect 93742 -908 192158 -868
rect 90360 -1098 141198 -1042
rect 90360 -1132 141132 -1098
rect 141166 -1132 141198 -1098
rect 90360 -1168 141198 -1132
rect 90360 -1178 90438 -1168
rect 85104 -1296 95784 -1290
rect 85104 -1300 106466 -1296
rect 85104 -1304 113234 -1300
rect 85104 -1324 115728 -1304
rect 85104 -1358 115659 -1324
rect 115693 -1358 115728 -1324
rect 85106 -1360 85168 -1358
rect 95730 -1364 115728 -1358
rect 106432 -1376 115728 -1364
rect 113208 -1384 115728 -1376
rect 81712 -1522 81778 -1502
rect 81712 -1528 87110 -1522
rect 92448 -1528 112832 -1522
rect 81712 -1532 112832 -1528
rect 81712 -1566 112794 -1532
rect 112828 -1566 112832 -1532
rect 81712 -1578 112832 -1566
rect 87080 -1584 92492 -1578
rect 78572 -1622 78754 -1620
rect 81746 -1622 81802 -1616
rect 90688 -1622 94746 -1620
rect 109150 -1622 109210 -1612
rect 78570 -1656 109158 -1622
rect 109192 -1656 109210 -1622
rect 78570 -1658 109210 -1656
rect 78570 -1660 90710 -1658
rect 109146 -1668 109210 -1658
rect 75524 -1714 105722 -1710
rect 75294 -1731 105722 -1714
rect 75294 -1750 105673 -1731
rect 75294 -1752 78622 -1750
rect 75294 -1766 75758 -1752
rect 105654 -1765 105673 -1750
rect 105707 -1765 105722 -1731
rect 105654 -1782 105722 -1765
rect 105654 -1788 105716 -1782
rect 75662 -1818 102084 -1814
rect 71804 -1832 71998 -1830
rect 75662 -1832 102432 -1818
rect 71804 -1839 102432 -1832
rect 71804 -1873 102385 -1839
rect 102419 -1873 102432 -1839
rect 71804 -1878 102432 -1873
rect 71946 -1882 102432 -1878
rect 75662 -1886 102432 -1882
rect 102054 -1890 102432 -1886
rect 68758 -1926 99390 -1920
rect 68758 -1956 99344 -1926
rect 68760 -1960 99344 -1956
rect 99378 -1960 99390 -1926
rect 68760 -1962 99390 -1960
rect 71944 -1966 99390 -1962
rect 99330 -1976 99388 -1966
<< viali >>
rect 97135 52542 97169 52576
rect 67662 52400 67696 52434
rect 96057 52412 96091 52446
rect 96285 52418 96319 52452
rect 97135 52288 97169 52322
rect 67664 51630 67698 51664
rect 93776 27537 93810 27571
rect 191891 27370 191925 27404
rect 198542 27392 198576 27426
rect 93774 27151 93808 27185
rect 191892 27003 191926 27037
rect 68764 48 68798 82
rect 115667 2404 115701 2438
rect 112790 1832 112824 1866
rect 109159 1671 109193 1705
rect 105690 1423 105724 1457
rect 102403 1197 102437 1231
rect 102403 931 102437 965
rect 105680 967 105714 1001
rect 109157 973 109191 1007
rect 102391 -679 102425 -645
rect 112794 934 112828 968
rect 141140 934 141174 968
rect 115667 864 115701 898
rect 99348 -798 99382 -764
rect 105683 -800 105717 -766
rect 112792 -694 112826 -660
rect 109156 -794 109190 -760
rect 115669 -758 115703 -724
rect 141132 -1132 141166 -1098
rect 115659 -1358 115693 -1324
rect 112794 -1566 112828 -1532
rect 109158 -1656 109192 -1622
rect 105673 -1765 105707 -1731
rect 102385 -1873 102419 -1839
rect 99344 -1960 99378 -1926
<< metal1 >>
rect 97118 52576 97186 52586
rect 97118 52542 97135 52576
rect 97169 52542 97186 52576
rect 97118 52528 97186 52542
rect 96280 52462 96342 52466
rect 96038 52452 96342 52462
rect 67656 52434 67710 52448
rect 67656 52400 67662 52434
rect 67696 52400 67710 52434
rect 96038 52446 96285 52452
rect 96038 52412 96057 52446
rect 96091 52418 96285 52446
rect 96319 52418 96342 52452
rect 96091 52412 96342 52418
rect 96038 52406 96342 52412
rect 96040 52402 96108 52406
rect 96280 52404 96342 52406
rect 67656 52392 67710 52400
rect 67658 51674 67700 52392
rect 97118 52328 97184 52528
rect 97118 52322 97186 52328
rect 97118 52288 97135 52322
rect 97169 52288 97186 52322
rect 97118 52270 97186 52288
rect 67650 51664 67710 51674
rect 67650 51630 67664 51664
rect 67698 51630 67710 51664
rect 67650 51616 67710 51630
rect 197006 27740 197116 27748
rect 197006 27688 197046 27740
rect 197098 27688 197116 27740
rect 197006 27680 197116 27688
rect 93750 27571 93834 27598
rect 93750 27537 93776 27571
rect 93810 27537 93834 27571
rect 93750 27185 93834 27537
rect 198528 27426 198610 27446
rect 93750 27151 93774 27185
rect 93808 27151 93834 27185
rect 93750 27132 93834 27151
rect 191880 27404 191938 27418
rect 191880 27370 191891 27404
rect 191925 27370 191938 27404
rect 198528 27392 198542 27426
rect 198576 27392 198610 27426
rect 198528 27374 198610 27392
rect 191880 27360 191938 27370
rect 191880 27050 191936 27360
rect 191880 27037 191938 27050
rect 191880 27003 191892 27037
rect 191926 27003 191938 27037
rect 191880 26992 191938 27003
rect 196282 26965 196372 27024
rect 196282 26913 196298 26965
rect 196350 26913 196372 26965
rect 196282 26886 196372 26913
rect 115634 2438 115722 2506
rect 115634 2404 115667 2438
rect 115701 2404 115722 2438
rect 112776 1870 112838 1874
rect 112776 1866 112840 1870
rect 112776 1832 112790 1866
rect 112824 1832 112840 1866
rect 112776 1826 112840 1832
rect 109150 1705 109200 1724
rect 109150 1671 109159 1705
rect 109193 1671 109200 1705
rect 105668 1457 105754 1500
rect 105668 1423 105690 1457
rect 105724 1423 105754 1457
rect 105668 1396 105754 1423
rect 68748 100 68816 1312
rect 102382 1231 102464 1260
rect 102382 1197 102403 1231
rect 102437 1197 102464 1231
rect 102382 965 102464 1197
rect 105668 1032 105710 1396
rect 102382 931 102403 965
rect 102437 931 102464 965
rect 105658 1001 105738 1032
rect 109150 1018 109200 1671
rect 105658 967 105680 1001
rect 105714 967 105738 1001
rect 105658 952 105738 967
rect 109148 1007 109200 1018
rect 109148 973 109157 1007
rect 109191 973 109200 1007
rect 109148 960 109200 973
rect 112776 968 112834 1826
rect 102382 896 102464 931
rect 112776 934 112794 968
rect 112828 934 112834 968
rect 112776 920 112834 934
rect 115634 898 115722 2404
rect 115634 864 115667 898
rect 115701 864 115722 898
rect 115634 828 115722 864
rect 141102 968 141204 1174
rect 141102 934 141140 968
rect 141174 934 141204 968
rect 68750 82 68816 100
rect 68750 48 68764 82
rect 68798 48 68816 82
rect 68750 28 68816 48
rect 102370 -645 102438 -606
rect 102370 -679 102391 -645
rect 102425 -679 102438 -645
rect 99328 -764 99392 -732
rect 99328 -798 99348 -764
rect 99382 -798 99392 -764
rect 99328 -1904 99392 -798
rect 102370 -1839 102438 -679
rect 112780 -660 112838 -630
rect 112780 -694 112792 -660
rect 112826 -694 112838 -660
rect 105670 -766 105740 -750
rect 105670 -800 105683 -766
rect 105717 -800 105740 -766
rect 105670 -814 105740 -800
rect 109148 -760 109200 -746
rect 109148 -794 109156 -760
rect 109190 -794 109200 -760
rect 109148 -800 109200 -794
rect 105672 -1714 105714 -814
rect 109148 -1612 109196 -800
rect 112780 -1532 112838 -694
rect 115626 -724 115726 -692
rect 115622 -758 115669 -724
rect 115703 -730 115726 -724
rect 115703 -758 115722 -730
rect 115622 -1324 115722 -758
rect 141102 -1030 141204 934
rect 141102 -1098 141198 -1030
rect 141102 -1132 141132 -1098
rect 141166 -1132 141198 -1098
rect 141102 -1164 141198 -1132
rect 115622 -1358 115659 -1324
rect 115693 -1358 115722 -1324
rect 115622 -1378 115722 -1358
rect 112780 -1566 112794 -1532
rect 112828 -1566 112838 -1532
rect 112780 -1580 112838 -1566
rect 109148 -1622 109210 -1612
rect 109148 -1640 109158 -1622
rect 109146 -1656 109158 -1640
rect 109192 -1656 109210 -1622
rect 109146 -1668 109210 -1656
rect 105660 -1720 105722 -1714
rect 105654 -1731 105722 -1720
rect 105654 -1765 105673 -1731
rect 105707 -1765 105722 -1731
rect 105654 -1782 105722 -1765
rect 105654 -1788 105716 -1782
rect 102370 -1873 102385 -1839
rect 102419 -1873 102438 -1839
rect 102370 -1890 102438 -1873
rect 99328 -1926 99390 -1904
rect 99328 -1946 99344 -1926
rect 99330 -1960 99344 -1946
rect 99378 -1960 99390 -1926
rect 99330 -1966 99390 -1960
rect 99330 -1976 99388 -1966
<< via1 >>
rect 197046 27688 197098 27740
rect 196298 26913 196350 26965
<< metal2 >>
rect 108964 51918 109086 51930
rect 108958 51882 109086 51918
rect 78606 51740 79736 51744
rect 108958 51742 109016 51882
rect 100608 51740 109016 51742
rect 78606 51700 109016 51740
rect 78606 51694 109000 51700
rect 78612 45584 78666 51694
rect 197030 27821 197120 27826
rect 197030 27765 197050 27821
rect 197106 27765 197120 27821
rect 197030 27740 197120 27765
rect 197030 27688 197046 27740
rect 197098 27688 197120 27740
rect 197030 27680 197120 27688
rect 191938 27330 194848 27334
rect 191938 27288 195816 27330
rect 194814 27286 195816 27288
rect 195754 26962 195816 27286
rect 196198 26965 196362 26984
rect 196198 26962 196298 26965
rect 195754 26913 196298 26962
rect 196350 26913 196362 26965
rect 195754 26886 196362 26913
rect 195754 26870 196232 26886
<< via2 >>
rect 197050 27765 197106 27821
<< metal3 >>
rect 197030 27915 197120 27940
rect 197030 27851 197049 27915
rect 197113 27851 197120 27915
rect 197030 27826 197120 27851
rect 197032 27821 197120 27826
rect 197032 27765 197050 27821
rect 197106 27765 197120 27821
rect 197032 27756 197120 27765
<< via3 >>
rect 197049 27851 197113 27915
<< metal4 >>
rect 98718 51758 100484 51828
rect 98720 51494 98806 51758
rect 98724 51396 98800 51494
rect 100396 51404 100476 51758
rect 76478 51204 82974 51206
rect 98724 51204 98796 51396
rect 76478 51134 98796 51204
rect 192840 29230 193268 29232
rect 196698 29230 197136 29242
rect 192840 29160 197140 29230
rect 196698 29156 197140 29160
rect 197044 27980 197140 29156
rect 197032 27958 197140 27980
rect 197032 27915 197128 27958
rect 197032 27851 197049 27915
rect 197113 27851 197128 27915
rect 197032 27834 197128 27851
use res250_layout  res250_layout_0
timestamp 1640022418
transform 1 0 67642 0 1 3396
box 218 -342 484 -90
use 8bitdac_layout  8bitdac_layout_0
timestamp 1640022418
transform 1 0 98026 0 1 1086
box 0 -1232 96520 51562
use 8bitdac_layout  8bitdac_layout_1
timestamp 1640022418
transform 1 0 0 0 1 1232
box 0 -1232 96520 51562
use switch_layout  switch_layout_0
timestamp 1640022418
transform 1 0 196132 0 1 26700
box 40 154 2460 1180
<< labels >>
rlabel locali s 198666 27404 198666 27404 4 out_v
rlabel metal4 s 197072 27958 197072 27958 4 vdd!
rlabel metal2 s 196242 26928 196242 26928 4 gnd!
rlabel locali s 198396 26794 198396 26794 4 x2_out_v
rlabel locali s 198392 27904 198392 27904 4 x1_out_v
rlabel locali s 196140 27266 196140 27266 4 d8
rlabel locali s 67886 3392 67886 3392 4 x1_vref5
rlabel locali s 68056 2954 68056 2954 4 x2_vref1
rlabel locali s 166012 3308 166012 3308 4 inp2
rlabel locali s 824 51932 824 51932 4 inp1
rlabel locali s 68780 -66 68780 -66 4 d0
rlabel locali s 90414 582 90414 582 4 d6
rlabel locali s 93764 2660 93764 2660 4 d7
rlabel locali s 85134 -908 85134 -908 4 d5
rlabel locali s 81746 -1340 81746 -1340 4 d4
rlabel locali s 78594 -484 78594 -484 4 d3
rlabel locali s 75332 -1538 75332 -1538 4 d2
rlabel locali s 71824 -1620 71824 -1620 4 d1
<< end >>
